�`���@^�T!�#WlRǑ R�������[�I� r{��|�������ޤ�#����$���~#5��Q�-dෙ�w�qIqR�T,ܘ�"�I7�!輫`�D48���I��φ��Í�2g8g_�WAv��=;�Hl�2�ˑ"-b9Vk����nߵ�9Y�B๮�-[��P������ǝ���i�\�_��k�	d��������<S�� ��cR�6 �o�1Y֎f�Xrޓ��E��H����1���i�F��$�	W3��dײG�[쏶�B��˹�<uJ˴��Y�TC�t�KqK�u�'ܙ�]/����������:���o��ve��H�9�Zd �F���Ȝ�Q׷A�Xk\aa^�=V���F|��KfC������rj:uÝ?z�
���ᝆ���5�g��V�XDf��z�|� ��Y�����*��,#׼_��RT�0���H���p����32κw�n�C�uu&�p�+7��ɢ�xa3�f7O�������]���wt1�><=s�;�H:��b��-q�(j�oN4�#�����8K�e�@��ƷX�Y��tvE{�����N)څz��-]�@�U��	_��v�!9�	�{�%C�Y����ڲ�$���.�[�~��>G�����
�9�n=ͯ�,c��"k�� f����H;�7��� G�����2�S�i�tqv:G1��:j�J�>t?��e�+���z�(��l�������Z�ףj�)�C�������σ#���r��(��SJ��a��Fd���n��5�*h���p����Y�Sǖi�/��~�����3B�y���1t�Mh�k�#z?�N�S��3��z�(x�6����8�F�����*�.���2|�G�~"_�鋌Tp��.�Þ�t�͉#K�Qr�\����nF����M�͂w�Л/z��%X�6��ϏM
�:���ġE���Q��g,%���=/d�3Í-��\�֢�@�:x������H.=�[N�בu�s`��p���0$�^C$�?AFEq������k�W!Gd��.�_��$d��d�Y6�mg�	~�'��Nb�x.�U���aV�Z�Aʞ�J�l��hh�i�B�r����n����/ܱ�o�W\��W���oH���I��=��BE�u��)A=�b=�ES�qpC��W�-��<�7�א���\�����f.�C!�A�$2Q1��Y�\g�2o�?��9��[ݑ�GYӭ�����2�r�Ўȯ�����P��R�1*h��#��h��m�p����)������]�Y�p�Z~pN���IJ�*��s�/=DO�k�}L�Q�Z������,��1�mwxu��Vk���:��N����|l�tV@���Z�fs�|#��i�'�mT1��Q[�1�]ݡ����8�Tyg��/xt�ެ����*~}䗈����@�,�6Hw�O�&�qބ\|�'M����`(�nd�d"�( �h-����ژ�-�Kc����eŇK��Xc�v/;�#���p/9Y��38�$8�|�<'��2�J�{(���&�J��?(�G}2_ �CK���cN��}#%��=� �>s��c�5R�����X�UZA�A;��R�E���MkKKK5%�V����c��}���ȹ�|����f�̴�"�$k���zj�4��O�h쫼qHX�]O�W�K�$��x�?O?1@�n,U���A���.�T:���#ݒ|����K����lM$CI&9G��i{���-�3͵��O��%�7��3�$g%�S٭�&��D�5y� ��W�#��K�~�+�hq���/����8[�^Y�g�1�6���?`�;��磚|~:F�Z�/>��u�U���p޿��%c�<��VT�j:�1��J3�<��aY�����T<�q~#�M����D�k�9;]O�W�f
C��U�tq.R�Q�7�+���b4���'F�jg4���4����qܠ_���֟�F[c&e0��;����f�!<�8�%��8P���q@�R�+�t���Y ("�ɲ�A�,U)'�*U���ԯՇ���P������)-W{��I�0���N�<@���P����7�c����k�#|M����h��C߿��ѧ3�%��P����L'�1��p�-�9wD��B�J.��E��b|:
1�t>:�k�=�G[���/�<Z]�[�wP�hoDA
���4�ʠͺx�p�9Թ�<c�H���)�2��G���6�<�B{�}Ѿ�Q�ϝ��Rnm�������.��=T��=�F��?��x��<��̱����-�U&(	p�����j%�R^7�u,(n��V��i��T�6�m�F#BIsE��udIF݇~&��#��aN�?.�?�#�� 7?�����Z�F;�G�����A�&jG�zD$��ߤN�����,5��!%7E�n������av��Uu�Q��9N������⚙'��"�=��TR��9EjZ>%�RV(g�6����C��}�=�:��j���L_��/�z����3dl3�?����f$�f���y���� O�E&��O�����e7�G!W���o:��>���l�Cv����򵤺p�3�%�����X>��=ĩ�q;���x�_Wj��x|�NU/�_����ޓ��P�H9]���-eI �6�ߒ�񥡴}���;�w�.x���^ﭯ�w���7�_@[e@9�������f�\����k�[=��Vl��eUlb�� ��3o� *���
���.��{�F��9�]T[�p�z]�[(&??o�~Rc��4i�tE�V��(�o���+O��˫��W�"J9Ņ3$+��[�jE���L��f��Գ�]�O�aߖA���>������P�l8�5�jZ@�'�g3�s�����D��Tq���*n��l�^���{�9����� Wr�r'!��c��SZ���j�t�C8��+4�O��X-ϋ���rOpL����B��RO���F�(���9��#����P�^��馞`��<���p�Hdȥv����D��M���5GtW��wO���(~|Mi��%�C���t�A��k���{�'�������m�}�u)?ӿ�VJk�5G"��B��Ӳ�A�%������4˼�,o�
��}B�>Fe��<#��j5�@�g7wG���G;�����!�8��V)��Vvt���}�η+;�4�(�qw'�v6���~�r���Ч)V�Cҍ�f���$i����M�6HiR:�x�tݐ	WΒ�K٨�)�?O�+ݗ�H_˿�o(U��J~_�e=����\)��R��5U��S�Q��<Y]�D�iݴd�����J�Ӵ;��6��~�R��h1ҍǆi�2Ș�&�q�%�O���陝cyݩ�vt��c����k��'�����K\%�e��6��/I����Grd$I�Ps�����j��/ZI��R�ʴ%�A��/�ZZ'HK��	�(��F+P�L#��ԸG-mVG������V[���v����	:\Ʃ�]}<���2ܝ�oΨ��*݅��9�Qsѻ�n����H�QaK��O�������\�7���~|'^	5@��.�JH�����ݟR�Lq��꾳>P��o��~��6T��1ܘ����j���cV����޶�疀
���p�:�H���l'��d��s��Q�(��	�����@q9R�p÷�Z��_bq��(5�$ɖ¥�������)W���Գ�c8��+�7|J׍O�:#��HX��v�8��w�0�g�2���Sb���r}�����A��T8�� �Ih&�5���%P�'�� ͘��+�I��҄�B�������V,���)�Q1���XB
�J���?r��L�Q˪��Y����*�m��}�%�icځv�;tR��}uI�F��D���IC1��ﭿ-d�����*NG8�<g�������Y���:��8�`w�{�;ߝ_�3�P�$��y�oM��4V���{(����c�Up�JK5]�T����(�.T�֣��~���?�U�Ψ�5�.��<s���z�au�y�w���	B��@ݚI���a�\NP
VM4	���4���:zc���W�3���o���0����9��m�6sM���H�!P��H˽P����Y`� Λs�O���-�h�N��mR���G��Eug+��\5Uۣ���������`H}�o�3�N{Ѿ�:���M�"L���d���-��S��>Շ��?@�/5V[�=_w��F����9�Wt���>g7泷��8th��+�'N��ϓ>�*���$U��ɲ<HΗK(ە@$�	jS�#�V�?�Nr��"�6=��4	�QŔ͆��I�/VK{�g*���Z��6\o��.Dl%�D�?�L�����x�[���S{�G�ww�RZUm�]I��h�4��Wv2����͇VM�����n��٭����4�3����lr�{�X���e���@q��!�,FH;�w�QH�m���xe7��Ju�zH�}��E�UB� �f����V՛�z}x����e�3��&j�C�3D��z�^�?r��f��|Ŀ��&�J����W�*�z,�Bi��JP�/�f)��5�J��+8�񵍪b��I�'��p�G����.����B��C�	(���Y�,�onF�M�vP䭎'&�����G|+�F#�����DE����}���J�v$��${�urEl�jt1���͇fm˵�Z���7��	ï��F������/B�KW��hxi�<V^!@ŔG�c����n��-m��-�0���)P�gx��������	�n��M�g]̅�@˲+9#�驞$oOu���p�m �" �Y��ϔ/����p����x5Q�R}���_--�k'�H�6RZ.�'&}�������Wi.eg�M��?<�����JF���<����g]��=��oك�'���;���u&8���r�G�]��nqϸ_��S�
�e�"6	�� q���_��ݖz`�/�W���J�����<Yݦ�Jk��J�� 7���D"Fe ho�EN��+��F����lt�z}�>��}��\o��%����n]A5kHث�/Dc^L*��_�[��V,7 y캪�XR�K�a�}����g�)�Fi��Qʌ1߷�YK��S��L�mˉv���� '���|�)����	�G?i�4L5N�J	Co��,�Yt���&���T@_s��fs��N�S��Ƹ�{�����sEx�"!Eh���z ��Lހ�^Zєp���-��R�������f��<��@&����F�%őbNѢz����,u������`�������O��ۘ���6GY�L�����Vo[;����q��W��
C@�{��b%������?*f�WP���c�=)o�'��2OY�TP;������W��{�I�zm-I#�	�!S�h`c���#��ùߟ�r��];�9�LB&���<ၷ<bq��@Y*R�.�=v��'�rYEF�TUO���U��삞5�;��{zy$��F�������E��z����{�uƺg����k��c�#��S���N9yO��xj�,#���w��-(�xq-��7���C�+o�x}/�@b�e�K��j{h�~�����j��ZғA.���I��޴?�w�E�����c�kU�jZl7Owk�5�:�hw�?�/��m�i�v�9����lxtm��
[��w��]�H��g�ϩ���g�wjy���T;����1�I8�FΑ�!(�O�Ģ�8-Eߤ�ieZ�֤uh}ڈ6��A�����s�L����N�'��'>D�/җ�+�����f}��Sߣ�c�%�.�Y��-����މ�v�v���k���R�ny��[ͭ��q뻍ܦH��k��ۂ��;�����gi�����О�@�]i8R�Xi<�i���4_Z
_!���H���6i�d�Ml�g�{����T�WkD���_�W�Ҡ:��VF���*\��5�JFu��k*Q��wہ7q����;��k{�2Y�!;�����H㤍� #�r3%1X]��hU����m�_ZCpYOx�R���U�5@�hCڄ�T�:�isښ���w�=P%o�N�at$C�щt*�Ngӹt]L�ӏ�*��F�.���Qz�~�TzDu�~�I�?�_���1-j���Q�9]~aT�[k��P��Q[�;S�gNw����˾��͙��PWP�n ��B��V8!\�ˊ����3r��\��Qׂk��5��Zo��'�\q�~^O@�zb�4���ϙw͝���{����LQ��{0���pRx*Fbd�R�0M�&��Zv�MBj��G[�u&K�)2���	�r(�=S���)��w�$j�����e�6W���E,?�2�hk&ߓ��.��wʃK�\Otm>��A� Ht?"�ՖB%M�*A^~S�rWy��C>!/R>W�Wd�s�@��6E������+�@~�W�=�/vA�[���>f�I�f?s0�h,�{�y����ɼcMt>t=1�=�a��L����>�I�'ɳ�#?S�񻓞�aZ���kP�z]tH�z:إ6���M����tGJ	r��#y�S�Յ�r�2?��F�~Zm��l&G��ć��t�o�4Kڮ��݆����|������Ǌ�e�~��Y�*[�||OZe>'n/G����b�3��}{���D��/B�N����;�s�%5NvG�U}�>W�i%��ʹH���F-C;��վҊ�&���7��Û=�{@��ޥ#�"d�H�@��)�b�be_�Զ[ڛl��%��:���٣Յ:�`a�0I��x\�!��R���N�����~9O~*WQ�+K����������j��s�`S�74��