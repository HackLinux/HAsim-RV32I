                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                RIFF�}  WAVEfmt      "V  "V    data�}  }}~~~}}}�������������}}~~��������~}���������}~�������~~}����������~~�������~~}������������}~~�������~~���������}~~���������~~}���������~�����~~~}}��������������||||�{�������������}~~~~~}���������������}}~~����~���������}}~���������~~����~~~~~�����~��������~~}}|���������������}}}}}}|����������������}~~~~}���������|�||�}}�~~�x�x��p��w~�~~��~��v��}�}}�}}�}��}��}����~~~~~~~�~~�}�}}���������{�����������}}}}}}}}������������||���~~������y~~�����������|}�~����~���������}~~�������||�{�����������}}~~~~~~}}����������{������}~~~������~~~~~~~����������y�y~������z����������~xxx~~������������u|{{{{�������~��qy�y��������{{zz��������xxx~�����������u�|}�}������||����z�������~�~�x~~~}������������~�~~~~~}}||����������|}~~~xx��~�������z���{�����|���������{��{����|��}�}}�|�u�|������������xx���yq����������|||uu||���������~~~~~~~~~~~~~~~��������|||{|���������xx�����~����|�{����{�|||��~~�����~~~~~}}}}}���|�����������}}~~xx��y�����������yy}}}}}~~�������{�}}�t|������~}}|||}~��������~~~~~}|�����~~}}x~~����������zzrzzyyy������������}|ut{zz~~~~������������}uuut{������������������}~�xyyyx����������||{{||}~|}������}}}||sr������������{��|uv}w~�����������xw~}|{~����}~{|}������������xwvmtz~������������zstltttt{�����������}vvvvv~~~���������|�����}~~~}����~~��������y�~~}}}|||�������~~~�~~}}}|���{���{�|}~����������xxwvutzy~������������|unogov~�����������zrrrrz�����������|unnnon~����������zmddldmvx�����������xgX[^jnyu���������zurwkplxsu~��������~yuunppwx�����������voh`^[]fq�����������xp\SLJNPbi�����������~m^WQMPThm������������ysnrnkqqrny~}����������������vmfceigoquz�����������tnbYQLHCCTl����������b216<@ABA?@U����������{E'&')+*1:X������о��lL;2-.5ALh~����ǿ����sfI@=AK[p����������k^XXXQS\g����������{_MHLQV[clt���������}raJ=236Kb�����ýï���uhYQDBHUcz������������tssy|~}wqj[UPSUoy��������҅<4;EJJKMLGG[�������ƿ�~G9D@?*%6l����������yOB:544,18R������������dJ?@CKU_er�����������nb`_o����~ssy����omjpv�����������ux}||}hbccr{������������{�z{qhdepu{{~|z������������zqkd\\_dcbj{��������}\Y]krsnllfbden��������ooy����qMFCN]l��������������zpc_Ycgq{��|y~�����������wsoljhhnopwy���������}}}ttsjriiiiy���������������}qijjsu}�������������~{y{y{zuuvwyvy|�����������y~{wtpmrtsv}�������rfqt������saWav�����wrgov������oc^fn~����~sot~������vrtvr{�����yzzzy�������yx�������{uw�������{zy�������{t{|����������||{{{{�|��~�y���������{z~}|{{�}yz|����������w}syvzxuxz�������~ea]p������x`]h|�����xmlqv�����ladgx������swz�����uvtwu}�����}wxx�������xzxvz����{x�}y�������~tz�~���|||}~������������~}||{�����|}~~��������~}|{{{{|}�����������}{x|ywtwy������|k_co������rj`d�����}piny������{peisu�����{wzu|�����qsuyy~������|uu{������}xurs�����|��������ypn|z~�����}|{����������{}wy�z�zz�x~���������~}}}yz{|xz|~������������{uzwywusw}������|adhs������pg]g������|onrz������uifjm}�����}ytw~����~~wytx}~�����}pry�������|wrwz���~�|yy~������yrxv|�����|�}z������|x~tyv�~����y~��������zwutt~x{�~����������zvztwxyxvx|�������vlcao}����~phegx�����ummry������ypflrv�����{wsv�������~|ttvr|�����|xtwy�������~y{vz���}vwz}�������|wyzz�����z{{z}�����}�{x}���|�z{{z������~|wyv{z����|��}�������|{yvztyy�����|onfk}�����kflk�����ymopx~����{slpmz����}vusyu�������wut{u}����}zvy|w������|yuz}~��~vu}~�������|wys||������{{{~�����}v��~�}xx�������zzvzw~~���~�������zzywswr}~~������ukhlu�����lgcqx�����{ojmu}�����uocgz������rqpv|������~wvuyy����}�tvy�������wuz|����zzvz{}������ylv