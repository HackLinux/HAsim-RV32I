    ,@MTPC7-'
 '*+/.)&#!!"!   ! 	          ):EOJB4*#
 '()*,)#            $0:C@82+

%+*&%#            (01-(!	 #(,(! 


	               %*'$ 	
                
$).,(!!                     #)22/%$% (,,)$	                        	%)431,+,( '45;6.'                          
"'.1656431+'!!##%(/6:>?7*                           	%,01469865520-'$%*019AB;*                        
%,046;A?>=;;91+%##%&+3=>5'                          )126768ACGA?;3-'"!.43*                            !'15:;41<<?A82)"
 $$
                               #,03-((026-&                                     #$#"$                                             
	                                                                                                                                                                                                                                                                                                                                                      ����    @   @                                                                                                                                                                                                                                                                                 
                               

      !&*&"&/5;:5.'    		                       	 ,8DJFB??ALPTTUKB8,  

                    "# '/;H\ntm_XWUVX[\`WRMF9'
	                    $*3;><;<FLUkz���zkdZYWVUUSUUNK?0                   
 )3=GSXX\\`it�����zslc\VOECCLUPIH>+	                   +6CMZdjpwzy������|smic_QIDEEJRPNC?1"                    '5AP]gpv���������xsieb_ZTPKMLOUNHD@4*                    
):J[jqy�������{uwpkea\ZWUSRRTXZQNLI?2'                   .>Rcqy��������ysqmgc_ZWRRQQSW[^YTQLH>2'                 #2DViv���������xrmhd`]XUROMMPSW[ZWXRMJ?5)                 $3DZnx���������wqkfb^XTSNMKKLPV[[XVTSOIB50&               $5EZlz���������yoie`[VTROOLLMPX\^\WTTVVOF<5'              	$2ARfw���������xqjc`]XTSQQONOT^efcZVVZ[XQJ?3'             
".<JZjx��������}vled_[[YYWVTW\fmojd^YY\\XNF<1            !.:EQ\fsz|������zrmhgcdedccbciovzunc\YZYWRH@2$            !+7BJRXagkty~���yttroooqtvquvx}��wmcXWVQLD<2"            "+5@EJNQX^ciq{�����||~~�����������vk\TOKF@6-            "+3;=BEHMRVZdpy��������������������}qeXJA=9/$            	#*059<?BFJLMR^ht��������������������zpaM=2-&           $,2457:=?EDCAFP\kr{�����������������ylQ9-'"          $*13457:==@<956:CMXgt�����������������~oS8*$	        #,247769;=>=830+-5>IS\itz~�������������zkV:)        )499<<;=<>?83.*'*.5>HQYeptz�����������vhQ7'       
",:>>?>?@>@>61+&'*-59BIPYelv~�������~zyuh\H8(
      $1<?BCBBCB?:4.)%(+.39=FKQ]gqz||��}~{snicXM?3+#
    &4?EEDCCEC?81+'&*-/354:EP]ehpolpskmoha\TIB<3/*
    *:FHJIFEEC;5-(')-./1/.5=KXadjhc`b[Z^ZSQJG>920-!!   -=GPRLHGGB<2+((+..-/*)09ET[\`^XWTNMNNIEB@=8431*#%(%	  	 .?MYZVPLFA;2+((*,+'&##.7BPUWXYXUPMIDB?<::;<510+!&++'	 	.@QaebYRIC:2,'''%$  +5EMRSTVYVOGA;79678:=50-)'(-,(
  ,?Sdone[OD92*&#" '5@LONPQXVOF92.0578:=3-()((,+(!
  '<Qfuxti[I8/' !###")2=HLLNQXWP@5,+.68;982*&'%(-2,&  
!5MastaN:+#"#&(*-2:CJNNQUTK<.,/269983,&"%',010(   -G]r�{iS;+$%&,/16=EKNMPPMC5.*./2682,'$$&(.785,   
'AZk{}xjW;+!$&(/37;DLQSRPNE:.)+,.042-%$$%&-6=<8.# 