GGHG�L�H��GM���������H��M���jM�jG�G>G>GB>>>>5>-/>=-57-C-===5.===?5??=@?>A@C@=@=\@?=D===5==5=/==--5=/=/>5B/>>G>>G>GjGGHL��H����M���M���M�Mj�ML��LHG�kk�H�����������������GjjGL���Lk������M�M���M������M���k���H��MGGGFG@E@>>>/--//-(---(---(((&&(PPOOOQOQRUQUUUcUccxzzz�|�����ււ{{yyccVUVUORRPPPP"#"+



�������������������������?=DBC@?BDDB?@@==5=?5-7-2-.-.(,&*(+(&*&+&&'(&&&(((((((&&*-&-(------E/E/>>>GGGGGGGGHGGMLML�LM��H��LM�LMGLG>GGGGGG>G>>GG>G>GIEG>�=.I/I>K���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I=@=���������&&&&(&&E--E>>>EGGGGM�M��M��kM�kM��M�|zxz}y}l}u&
-(((-&(E(/>>E>>>>E>GEGGGEGGGEGGGGGGHGGGFGG>FGGGGGEGG>E@EGGGGGGGGGLHGGM����M��M�k��M�M��k�MkMjH��MjHGGGGE>FGEIEG>>>E>>/EG@GGGGGGGFGGHLMj�����k�H�����������HG�G�G�GGG@F@>/>>@>5/=//--7/5==?====?=5=BCD@C@BCBA?=B?@?B?=====-7=====/=5///5>>>>GG@GBGGGG�M���M��k���M����k���H�GHjM�LM��kH�����������������GjL�jL�HLL�M�����������M��������M�M��H���LHGGGGE>>>>>/E-/--(--&E&--((((-POOPQOQQQQUSSUUccccxz{|{��{��|||{{xxccScVSQRQRPRPP"""-%


�������������������������==CDCB@?D==BCB?==5=5.(5,-,-,*-,(*(%&%(,&%&*&&&&(((((&(&(*&(---/--//-/E>>>>G>GEGGGGGGM�LMLM��GGMGMLHLLHGG>G>EGGG@GG>I>>>>>>IE%�?(=@?IL���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I=@@���������&&&&&&(E&-E>>EGGGGGHLM�����M�kM�M�k���zx{y}y}uu&-(-(-(E&-E>>E>@EG>>GGGGGGGEGGEGGGGGLGGH@GHGGGGHGGG>GEGEGGEGGMGGHLH��M�����M���k���M������M��M�M��j�GLGGEG>>>E>G>E>>GEGE>>GGG>GGLGGHLG����M����M������k�M�kL�MGHL�jGLGBG>>@>B>@/5=5/.-=/2?>==?=?B=@?BJB\@C@@?>AD=?BDCB?=>===5=@=>5=/>5//>/>BGGGGIGjLLH�����M��Mk��kM�����M�M�����j�k�kH�����������������G�j��j�L�G��jM��������������������H�MLMj��GLGGGF>GE@>>--E--(--(---------PPROQQRUQSSSSUcUcccx{{||{|z��|�{{zcccUUUSUQQOPRP"P"#",&%

�������������������������,=@CDDCBD@=DB?=B=5=.-,-,,(,-2(,*(,*&)&('&&(%&&&&((((((((-&-----/->-E-//E>>GGGGGGGGGMGML��GMLMGGGGGGMGLGGGGG>GIGG@G>G>>>>>>>>&�@(@I=IG���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.I/���������&&&&&&-&--E>G>GGGGML�M���M�kM��MH��M�|z{{}y}u~u(-((-(-&E/>>>GE@GFGGGGGMGGGGGGGGFGHLMLLHGLGHGGGGMGGFGGGGGEGGLMLML��k��M������M�M�������������M����MLHG>GEG>E>G>G>G>>>>GEGG>�GGFGGGGHGM�����������������M��k�jLGML�jLGG@GB>>>=B>=/-5-=5./=?B?@=B@CBC@\@\@DBCB?@BA>C@KBC?==?===>5?=5=/>5>5>/G@jGLGL��H�����k�M�M���M�����������M�����k�������������������GjG�LL�G�H����������������������k�M�k�GM��M�GGGGG>>G/>>/------(---E//---RPRRRRRRURUUUdVylxyx{{{|{|{{|zzzzyxccUUUU`VR`PPPPPP"P-&&�������������������������,5?\D@D@CD@@=D==?5=5,-2-,*(-.-,(,(,&(&+&&)&&&&&&&&((((-((-(--(-/-/---E//E>GGGGIGGGHLGHGMLLHGGGMGGGGLMIGGGGGGGEG>G>>G/>E@>>/>&%�?(/@@IG���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.?>���������&&&&&((--E>G>GGGHG�MLk��M�Mk�HMLH�M��{{y�yuyuu(((-(E&E-E@IEGGGIGGGEGGLLGGFGGLGGHLM�jHLLHLGGGGGLGGE>>>GEGGLH�H���M���k�M��M�k���M������������M�k���GGEG>GE>>GGG>G>>GG>G>GGGGGG>GGHGH�������������������H�L�HG�LH�LLGGGGB@>>/B/5/--.5-75?=DB?B@DC@D?DD\BD@=?BC=@C@B\@@?B?@=?5====/5-//>5/BG>�LGG�L�����M����M�k��M������������LMj���kk�����������������GjGj�LjG�G�H��������������������M�H�M�H����GjLGGG@>>>>/E-(---(----E///E/RQRRRRVVVVUdUddyxdxx{{yz{{{|�{�{y{yydUUVVR`RRRRPP"P""5&(&%�������������������������,5=D\@CZ@DCB?=>=?=-,-*-,(,,*=2(*,(*(,%&&%&&%&&&&&&&--&(((-(-((-------(EE-/>>GGGGGGGGGGGGGMGGGGFGGEGGGHLGGGGGGI>>G>G>>/>/>>/>>(�>(@?@@I���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I,@>���������&&&&((-E-EG>>HGLLHLLM���M�HLHMH�MjM�{{yyy}uuu(-((((-(-->EG>>GEM@GGGGGHGGGGGFHGGHL��GjMLMjLHGGLHGGGEGEG>GGHLMLj�M���M�������M�k����������������M�k�GGGE>GE>G>GG>EG>G@GF>GGGHGGGGGGG��M����������M�����k��H�G�H�L�jGGLGG