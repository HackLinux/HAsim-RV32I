{��.jK�p,gN�H�Ii����ܰ1R��4���*���C�-����/jL��������T\ޝ�|~��-o��k�nʝ��|α�8�!Kv�{���)Қ����dr&+\��q�Q��WϚQN���7�Db��Q^<�En�#��V9�II�x�i�c�-��|���ߖ��uD��]�#{+�3�~!D,�e���F�f���q���X&L�M��S?�`��x6�]�M�"k�ǭ�Zױȯ���Uc��MP���!IV[1*ǔZ���GsT�s�$���>� �1�~�K�\�����D�/���s+�Ҙ7�S2�T�_l A/]W^3)}�Z����x��ך0�m�GE��G|YrEo;EA��B<���E��.�[k����py�,}��KQG�����vĮr�mՑ6��
^��~hh�<�b
���?`�Əǌ��a��v�D�[�>g�S�>�܈�H�?��7Wۏ&�i��v0�$���d�槪*�*ѯ��w��"s#�T��tZ���m����ܰ�S!��;�a�lᴳ���$�W�n���q(���UT��h!&NT$�6/C{��d�2/�IT?oG� |"����4)m��<����$���S�uҺ����4���&B�CF�W��� @6��z׶¨���9�Ӫ��qŭ���&��o�yF�,lt<#C����9�ס����kq&����as�������V߁�>wa�y�p��ǡ�گj>OoZ��s�fh��_��3�t��cJD��Kھ<̻`�L {��a2�ѳE�὏m����l5�!-#��n�d3�i�i��ʁ��ژ�P%H��� �-����Ղ4|���KIѨ�ШOV�[���&Q�]�@�%G��v�'oӪP�����0����N掠����l<���@��y��n�1��VM�]. �vz�6�,�-��t�E5Q��q��
Pr ��1Xd��<m'T�pj&�wk!��vl ��qm'T��ﮊ��lP����h�	J[	:
��~&�}�sA��Z���z�-�;��[g�{`����t���6g���'�8z�iI�c:ZB"��|:�f�������V9�����o�fW��q�|sZH��o� 0�����7.xF���x>�GwʘJz�ʜ=t�:��3����wv ��;ש-�g�:��c�T}�Q�UP����� ���@������P�T�ڲ9_B46��j+�|�Q2®�0G���y�?B�UI[7����uK pP����E�"{CΈ�e$q G%YȴI�t�������өi��nv"��'UaJGX�uȊ,�N,ӿ��AKDQ��GF�euRp��!`gj٨b�z��Ӈ1�â~��g��%Vv���tKq���jc$�e����"]���l�s�B�(�������a��!e52FpGB}rp՛��1��p<�%�S���tI�a�*�yeR�?��V��ic���H�$@�ǘ���~��E��d�-bg����̴cD��`�٠˴K��++"#ϣ�d:Y���3~�՝r�j��o ���h�Ċ菢u��A/�d�$$�o�����҉����=L�:Ŀ�R��ӤK�����m+��D��5��Q��K*���[����rr���"���**3�fbo�g�.��̈�+���7�_D�����Rf�""�B�/n��Z�ٝ�c���hƷ�R����(���M���C�#0�@�1dL8�W�v��3���:I_�q��e����{����@��QQ�J9=o�p:�f����P����*X/�k����wk3�X������Xz:n�సT��{g�������]�zp�.�S:4ΒWcѻd�%#��,X���H<OO^Q�,�*���	�y�fu#A�8.��b��wft��~At$2!Ƶ�cJY7v	�/M�����<�dU�Vù�:��G�A��.�b����G��MuB�����x�0�j9��4Y�4�3j�Rk-�S��?x#��.�h\�ӣD��oԄA٫��Y���e�K��m���Qk�>�0J7I�eы�Q9�O�)_�tD�@�1����Scq���|��� �# Zv��Y �Pƃ��4�ʗ�I�ƥ1�9XG�}܆���:�t����ɯ�R(�b�f� �P�u������t��IJ���	r����-i�i>����L
��b�`)X���+��<Я�l�l���ǵF�Bs9u����e��jeQ7p��Δ,Ë�4�g]�6Υ��]���q4���F%r�g� ���q;�nO��lǰ�T����q#(�t�~u�A�G�z�x�pž����ٟ�!�h�/\5���,�s6�A�]�9R�W&�9`���!��S����iғ�iGd���G\ q`F���|� �oU��D`ۻ�_sf��O�׌�W��Q[�n���S��.y[&�e/RK1�
5��a��A{�\X֜����_0�|��)��!��bf�YwMn;�i�Sd�� yx��my����|�9��;*�9E��W�K5��k_1�æQ���afgC�z4���8Ȃ�a�uZ��2dۏR�):��+�j囯q0>����GRv����c�˺v� Q �@��E(3�`�8��B��x2��b��4Ij�	~��J����Pž~�q��M�~�v�9���^�_~74�I]�H��1,JpT�$w���e>�����¯���C*�9X
3D��̮A���,y�Z�xmAfLa��o_P$�@�!;ç-6 k�)2��#�(iB/4�!�/E���"�n��ʁ��}�a������P%r(���(L�7n��$�y�����n[��10���w���B�B��;�4�m���v�2������ە׏;�Q�̨GD��eۥ^�֏ܣP]�s �����dFv�ǯ엺j5E��v=ViƮ�V\���o�E��ۂh��*Ax�KE�.gg#LOT��t�F1ּ�q�-c92L����� &Bv�G�0k% w���O�x��K�$��˴:�U闘MpN�9�,�N�V��S�����5����Va�=�Х��?����ofG�4�|��}c�+d�ћ&��n��<���'t��ӋE�z� ҒťC�f�-��8g������$y�����r�G�FW>F �D�>t���F��:���������
�tk����L�*�R�f�Y,�.�	����2�'����H�m3�1D�<~1�M�L�9۹$~��F�ƅ����
 ���x0[�d�T��w�E�-4�H��� 5��!����X���ըr ,���b�)CO�D��!�b�TMΫ��)��y7o@i��>}��D�7�˽�%��feC��~���FpMX �2���x4X�o�l���p
Y2�O>hd"l:��K��N���sĵ�����V��8>���AIe�3�v&�cY��oE���L��<���k�Y��<g��yn��)�tZMEw�ʌ��>8yt���K�9!�|�yB��E���ǌ=`�U�܉.�sm��?��A�����ܡen
O2��Vb��u=?-����B�� �jۂ5v&/S	#�6��C����\�
?fOv�W�΂OX ���k3=s�p}\z�Ժ^G��o�M�#�Y��PG���>�^�{�^��0
�[��1O�9j]���l�/���C����z�I��c�	Z�bӇ�I�H]���	
s'����F�����/�~� ���v��l�NԼ����b�30{��~ӽ�0ї�q�p-����f'���z�A)��~6^�!�0 qq�!n�����&%��k�]w���A��Q������;z�N�M^�Dk}�g�vY�A���UF�a.����싿M�+5�r��_G�)6hM5^4�7��lH��`�hL�M$��,�K� �-5G��.t�H�Nj�2)��;�a�I��(��0����z)�p[�3N�o�,٘Jv�ޝ�j�)�҈nʳ>kU�wa$��&x�u�N�%����A�>{�a�-S��j��?v�jL�W�1�+�H�4��V˥p�=9�_�V��)�9�s��|W��|&��C���zp;W�}l�c6��j-���|�+�D���$��fZ����{��*L����vF���$3�{���^��*6�<���Ï�k��o ���O���������L�aI0�uve��$*���S�������WI��[`��l<7�nGp�e��M_+ʅ?��]���t�A{�2@=������0R;B�r��