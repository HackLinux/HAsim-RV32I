UH>0 )����yvovz�����y�yjijnkcnji^jz��wwunvzjg^Uy���yvwwwz�����������jjjjjjn��wnj^i�����zyz���zojnonoy��wonovvwwonoow���������������uuvwz�vno���z�������wvvvonnji^i����zz�������������njouT@U_c]U^UE0G����vvonn��������jdiii_njiUcy��wvojn�wjgw��vjidjjnno�����w����jfjjfcn��vjfci����wvwno��������w���onkjjfidnw������������������vnoovwnio����������ywunnkjji_^fjo���w�������������vnvvQGUc^TSQL>)8v����wvoooo�������vj_ejownjUXwvw�vniiw�����_'';_nniv���������wijijio��okjgf���wuuojv�������ojj��onnkjj^U^j������������������ujnouvjivvjn������wwvonjjfji_jmjcv��vw��zyy�������wnvwjGGTPEGE>8Gv����wvuuovnu�������vjkw��vfiionv�wnidn����c'+4('"4]T8d����������njfjknwzonj_n���onkjn�������vjc_iowonnonjd]Tw�����������������vnonnn^dvvjiov����wvuooz���zvvojiw�zow�zwvqz������wjoyviLSGUjjjcn�����vovwwojjw������������zuovono�zojjn���w88HSG8'4>5,8gnnv������wvuoojnwonjiy��wnjjonjjo����njji^jwwoonnjj_Xw��������������ojzwnjjjjXXvvjjjdjw������������zyvnjy�wnv�wvono������ynovzwnoow��yq�������vvvvojjn������������yrwwvvw��unjk���n;GX^UG4@ADHE811_w����vvonkmvwwnjjf���vjfnvj^TG^y�znjjf_io�zunjji_j������������