�>�R���B
1J$�eu�(�ٰr��/���MQ���d�����S5�
AگA�|+�@�sŏDy5�&�nt"�v_�{E6�x�h�pAz������R9�P��1j��<=���r".��X��[�ri"0թ@G���!Y�����cs����#��V����)nC��8�F��s�F�cs�i;���T�\��Y�^ц0NŔS0�w�a�����9K\P�o�1�������AA���k'�>w��sŀ���͠	���T0��4�2�F��P0��4p���n��Z�G���ᬉE6�zo����`������nӂ&ct�����)��as�����|��s�^ֲ���4�A@%C���&�����p����eZ�2��z��.�x�4�zD��D塹����Uֻ7���5Er3�Цf�y�薒�7���G7ħl�����������#񶒋EĢÀs�������&�2$���h?���]�7���B1�Ѕuc�����yj����9�G 7慠��k̬uۇ3��?����F6��>AړAtu�f���h3o�(��t#�e�kk���δ������lc�����Ҫ3F#��t�߉t$h=�����A-1�%Cs�����@!�̙�e�Ar��PE��t�9��ۣQ�G7\�U@�Gۯ��nq�G?7\�A@͊��YF��Ǩa��w_�o�Qф��?�(`s@u��`���UЁf�@n��@�d�97l����y���J\��S��qF[g�������Jg��aEi&yO&�VэZCAfc���x�BB@a�Gu����t�7��ef n����Q��X�� p�,A"i��f��bE��_r���]֩F*E&63�{թ��*E6��t� G�Ǣ��rŨ���t�Q���d�L�,|�@gm�����T�1��"Rv�HGlxE��iz�~{K�bB���#�\�q�nK@�P����^��iҙ�$6�B�!�o��YЀL�/%�?�R�<�,D37\�?@5zx���7s�4`���`�`ʅ�$�ܣC70!��}���$��0��j0��ĬU@����y0Q�y�! 0��>0����_@��"��i,C0�+309=r�`A"�@s��f]���j�j���ab	�����V�jC'1��FS����s�ֻ~��&F#�Qt��1Z���p�鷆�mV�}� %�`��u+���j�}Z�!�o��?�gW�q�F�گ�y�W�9�U�{�V���i!t�97����re�/����襛���aH�s��<7�E7|�@E�'R�g�SW�g���<�T�p�gFk@��T�u����l��m�n@*@�E��b�􊔬U@�jr�CFS��Et���t��J��}Ƣ�uĭ��]Ѽj�B�`����Qc�3��o"P���^��&�Ʈ�֮�G�|uF�u���)�(ʩ�>�$1f�����4�ݹud��g����s�ѽ��9'CG�C�~˩���~�U�i+P��w$�q]�\h�u�'W���o��nѸ�E�����b�����ʎ���<A���PVf�D� ECG���V�I1������ͯ���o�l���w�e]׭��Y�f�� ��鐌���Agq�y7��6��R�*F����7�k �0W��� �#6&,A"`ې+G#6A�ʶu�Ft#3t����y����+@1
��t,������]V%�_�M\֝C-0-����[@���)ˮ�����$m���.��ˮ�k���Tp�XA�A��0s�z�]�����LT��-F.7��z�rc��]���l��b�]W�W�~�[��"��se��S�x�!mA��|������3.��`"�fa���*]��� 1��60p�e����˩t�,�˅�H.*@
1&W�f��� Å��{�g�$iJ�\����@v@���˹u����UP�o��j���ƨ}���n�a�e褣��qU��k`�K�)�A�J�䢯�h%ԁ���0���h�u��*�7��o���@EkG������������j&��:Tt�}@�����")���p�t�g클4#c��Zѯ�+���"�F�o��G��u�Tt�2����k+�����+cGdڀ�&��u����2A�bA:�~A:@��h(4��p����F� ��vrG�}I������7��S�����W�C���
�X�/7����r���b]P�����TuW���w�B�p4A2���Y�Ć�KS������A2n@0+�Q�X��re��u��s����6��d6��6toG77�o�7������������ ���|���&��LT�C'��Q�|��e�ك7��C,0�&�T�E6���6���l"����ƍY֏�����mS@���qF�!柶��pm+F레�n8|�|�R�1]Wj"̈��B 0�5�R@{��'h*�<1&%�%uÀ���⡤���{ECG����F�^���t��M�_�nѿ�L�P������(�I����!eA���C�܇E!E���41&����0���_��Z����R�V�v	�Su�u#�e����e�ٵ\�zX�4�b�T�h�s�y��\�Vѥ3�r��O�n����M� ��(�ҍ줊�K�f����� ��z�Wь[좯��F� �Ư��<ԍ�	B0}�*G�ʉ��d!A&BYse�_��b������u�}ũF���r�&����m〼��a���ϓ'J+Ŕˮ:Ar��juD��u�s	��������(�qx�o�{@����A�s� �켞@B@�N��y;�����'
0ez�����ʎ����MX�mB10�4�h�~�3���׃�6����	[P�$Dt��	t�H߫t�Юt������0~߯0B߬uD�qt�C�)��T-"��.q���g��1��mv�G��g�U���c������F��)s^aP���rjaP�{������#qՐ��a��iw��c���[et���2�	0�d��66��h��L��L�,g��7�(�r���.���B����G��\�j��g��d���
I��y_aC�����t�w�6�5�A��qu�ʖ�����Fb�u�"��gw�G|ƥ�X��v"t��9u�n�:����W���߳g*C1��v�A@Ac����LfQw�'�=�y-�V���im��+s�穀����;r���a�zUP�6���VD�x��G��<лx0���,�+7,�p�F#��X�e�$=6��-������ݩF�*ʝ��D&6�xhFkb����K
ʝ�}����/f����%�����<A��bt�v5�J��=���eu�����BUЬ!�vZ��������&�������r-��%���"���eA9Ajkw�~G B	054�#�~&v����&4F���i���W�*�����d3�g���)��a����x$���:FTF��xȮG�Ղ��׀�b��=xUFxz�a�^�o���ڮWy$�7t~�7z8���7r��H�i�8�M[֩���#:ޤE-7��@#1�|ʨ�� CvԮ'iN���0���,�G6sxϯ ��sEǽφuc��Oi���6m2��m'4Ӿu#��O��y�g��_Q�ḌP��"0=4�PA��r���(��O����|�0�[FC!��s��T֍D4�A���A0��4(6�c�Ϡ���&eC^�-afAz�1�G��4��"� �j��I�f�X��t���h��O1��2I�䩦rj���g�T� ���^u㩷Ɉs����S֡Mm`rB���p�c%C�H����hfE�/�n��I�m!���G�������P6����d0rb�|�1�a�J�Fg�ʇ�[�0�*G%ՠ-��&���6�&��QV�"#7dt3�iF��]ї#V���҅4)�(�`v�@m���̯�t�x��p�׍[��*F+6[A��vt�����Sך�w����fI`s�zA2�w����ЌY�������㦗�%��Ư�}�������Vа��6��a#��u���ы\��B��t�,y�����́����}��s���b�L��1���jAJa�¾t�-k�7���۫F@��r⸆q^�
C&1�B��
�w�q�����+�%6��JA��RA��BA���w���$����-�YГ�hF�*,12�c�dr"���i�z�����w��ޮ�&1j�+Fg��pL��8��Ԓ����{"�i�� ����drm���.���nq̖���s��:c���t�Ľ�8sg_���(��?�nQ��H�~�P�����xLY�������E7���ցt�K�.v�~)@�h��^�|E)7\��C'1ګoF���eu��*�Y���'�ӱu$�.����X�+~��{E�-�Ȯ��)��AA�M}U��&���s���7���!I}V���C�{��V׺�����hE07C|����W�o�&��P�r�+F� �пr�V����iFÇ�eu�`���ӱ��;�B	0�|��vJ�/�����#�%ex�gT◗g~̛�e�DG������-�T�[
�aͯ���̾yK\�����
�B�V%�6��B0����u��<�{ݩv��drbM4}����~�W�'�RQ�%6��y	�d�c}����+��0̿�ڶG�}"C"���[��xA7���7��77��� �E66��Z+N���v%��u�MZ�C��[��|�9��E ��7��{ΪA����������������T��1ʪq�J\���rbS�p���De�7}#1�@��׃��|dq@���Yu��^��5_֪$d3��t����dr�8ABk��Y֫�p,6�|DA�}o��r�.��x�cF�������@�?ZPoq�{F�+F{$��JV�wU�r���#��|����*��Lp��*�ڰ�D����A�@���ƫG�ޭʶ�]���F7���!���酣�or���)���A6��L0�~{�KF׸�߶��K��<�