%���Ȁܤ��.�-�"G!D̅������%N�4�TC�s�<xe!������%����Q�N�wib���%�a���u�^cwM���nd��%���$���S����"3�Q {`����U���m'�L��m]aN�J稣?D�f2�$��3��j��G�9Eɲ�)BHL�#C��[�!� E�/B���~9"Tk���u)"�ζ嫂�ܕpH��Е�0�ݕ��K��(����l5�k��k��݁�#��Vؕ��\���_dWf$Ne0�'#[3��J3�����(�N�e�c��Sԕ�_\��D"�ܼJX�ۏd���L>#7��L���Y1b�n�K�Aޓ�Z����ƒMX�Z�(dcF��ڽ��ߕ�I�siM'���$�N���Fj��٪$Jx>�޷>,�L��ǻv��c��d\c,r;4��-��Q�nM��I-n���CȪ*��wO�wl:?
XB|U,ڊ!�I��c�U�������)��_����4Ȉ�q��ICF:>��P���7����H0��ĥ��o�C%�b�$H��RVc�n������o;4�NS��N�Im��A������/�Ϙ�BG���,�K�îxw�N�l,0��.��	�U ������� ={�樌���-�N����5��2������dA\��.�X�Q�Sb'�B������n� CiyV���D�x�������姮��V�3����H��$��K�v���֫�g厪��dL~Χ�Ds����&O��u������c�n��G�35�q��n��G
����D�W�@ND�52�a���@Yb�U�e��vA�Jyj&fßj,��B��y���^�β���)��!��f���v��<��:l�U�2��lj���"���3���X��۠� ���}A��f���{�}_!s�n
4��EѮf�w���M���[��qt��*�6��w�8����,��$F�2���X�|2޼��_w�q��Y� � �I�����qƔI�h��濥#�8׌��j#��TڏU�0��d#��d#��<c~K��`�=zQ>�)-? V|�+�<9��Z����|��A/a��i����%W|,�����DO��o?��ء��.+��y�bX�*9:�uo/�*
�g���$�
�S�cF�oI)Zu֛��g�,�C� ֽƤ֭˫���{�N�{��QY�E�#��;���ƣ�ޮO�$�ՑR./��X°7�(R,(���3*Lq��`���jt��ء�;���m���4V�a���$ċ��&�/ ��81�Mm9�x� ��V5�E�~6�r)�4��,�2=
�v�Q�#Yu4����n��ńAA�L�Fe넓Ǽ�|36 �b!�y�󢖅d�F��4�z��3`��T`��x�
:�7CB������'����8��+�ɈK'�Vb����n!�d#T�q��h��Fxő�J�U�hV��;�5}ȱ��1�i��?�\��H�w~��n��8�RXsZ�E���G�[$p肤�j�]��b�(�n�Lo��b�,�f���AQ�+��<�]�������孮x]^�������*-���~�N��d	��`�