�3k���BNS$5�D A� E$�ND�N+�NC�T<�VB}Y?<\!t^�bD�e;�e=fg0+gBn.oA�s?�w6nx$��A�5R$S&�S�b�~ X�,'�$�e $NS-�],ag3kp
�~#$&�W%Y'c[\6�]8�e<eg0fk7�y"I{<�*��R�?h�:ň(�8Џ)Y�e1 @2 K$* N
NJN5NNDN]$NC*N&-N/:NA;NI>NQLNIYN]�NV�N8�NF�N@�NN�NP�ND�N@�NO�NE
OQOKMOX�OZ�OBDQ]ZQThQ9lQTqQYsQRvQNwQLxQ\�QG�RHS_SUASQWSNpSJ�Sc�SJ�S4�S6�SQ�SW�SKTP	T[TZTW&T(�TN�T[Ua/UE�U]�VU�V?WY(W0fWU�WU�XPYD'Y@)Y2eYM}YK�YG_[U�[G�[R�[U�[J\P<\Oq\9�]N�]=E^c�^O�^U:_WS_=�_]�_E�_L`IP`[�`YaVb7�bV�bQ	cWwcZ�cWidX?eV�eL�eP�eH�eO�eFzfR g/	g:gP*gX,gI�gU8hW9hO'k8dkYlT4lL}l^�lT�lU�lK�lP%mZwmL�oN�rJ1uC�vN�vD�xe<yZ>y@�ySFz`,{9�|]�~]�~J�~O�~O�~G�~9\U`WT�>�`�PT�<��Y��R�K��D6�U�Va�^��V�E��^׋^�J�U8�b^�T��T��Yя4ُ@u�`��O?�Jd�^��R^�@�M��A��Hl�O��Y�W�TN�M	N.�_"6q&v":y�dqfNf�bgn(�')R?NSB�S	T")Y-:_:�`4�g#�l*1m<!n>^tFW)��0	�@�M�@�@&�6S�6:S�_l�l(�p$')R�R�V,�^ ga�� �3��"N\P�e!�Q)n�6R�R�S��R�S7OS#[W.�h�v3z��,:N-wQ;�RY}Y"�[9^5�^,:_-�_2�e./f 	g(�m9�y?wz@�7 �0�y���Q0R>�T1�W1{_wm"T�17��N$TNENPNQ%NT:NE;NDO;OLNO?sO0�OPHQ<wQ6�QQRNSBWS?qS^�ST�S?�S?�SST4}TPZWX�WUYA'Y
}Y1�[]�[V�[@\I\V^M8^Vr^\t^:^5�^v:_F%`c'``�`3bQd`�e/�e$nf`	g6CgLpgTAmP�mUo[no]kpS�pPrX[rF�sVEuF�wT^ySwz[�|VA~L�~[�~<:Q�4�NP�eW�>�Cj�c�T+�F5�RZ�aя'�P �<v�Zؚ7�QN�7Q�OR�9� �N'�N6R,c[0�[8�[/E\1�]4�^4�e-�e/g48h=Gl-�m1t&u7��.��*^�*|�(1 <2 B3 G4 J5 L6 N7 S8 O9 VD e$0 N?	NQ
NZNRNfNTNj$NP*NM-NB0N];N_IN\]NofN`�Nb�N`�NU�N[�Nx�NN�Nd�NE�NT�Nj�N_OOnOaOOVSOjUOd�OZ�OXEQfhQ`kQglQMmQlqQasQ#tQg�Qp�QK�Qf�Qs�Q_�QT�Qd)RJ6RMoR`SASi;SUASWUS?`So�Sm�Sr�Sk�S8�SE�SK�SLTZTgTF�TE�Tl�TfFU.�Uq�V\�V_�Vc�VVW2:Wh�Wg�Wk�WgYnYKYM'Y)Yh}Y\�ZmX[Z_[v�[h�[W�[i�[l\o\:E\b`\mq\k�].�]g^h^g^Y�^f�^Rq_Q�_I�_N'`j�`\aTbabXbq?bXybW�bP�c69el?emHeRpeY�eV�ec�ep�eh�e^�fY	gkgrgP:gQCgIagZ�g>�hg�hV�k}�k|�kj�khl@4l^}ld�lUAmS+ovdqDgqpirbyrS�r7tguc5uV~vU�vG�v^�vZ�wZ�wO�yj�y_�y] zv�zf�znI{m�{p�|8�|j�~b�~J�~=�~K�~*�~p�~uDy�LK�xL�eT�l��_��9��L�X*�go�gr�<ׂnR�ao�`܃L,�W��`��GƋc�r"�M#�]8�jD���c��a��c��\Ǐ_ЏbяJُS܏p�YёM��l��^��g��B�o?�nP�Cv�pƖT��^^�j��f��lߘU�hm�mn�o��n��Uؚh�I�k�\(�[7�3N�:Q�eKQ>�S R;�R�[My_?�v;,{Gňp�&��ET�G^�e�f,���N3xQ<Љ#!�:Α	��7�"
R^7�_g&�v<'���N-�N=vPpQ36R+;R0_=,g-Pg�i4Gr*Hr0u6��6�'Ֆ-�)�S:1\Abeg�k@>m4�~0�~A�� ��=�Nt^g$:N%hT1�V*W	J\6�]Et^0�^@�b"g&eg+�hL!k@0uB�y2I�9"�;���/��F�(7�(;` ���q $�S�b!kO4sQ16R?�R,hV&:W �[E�^$�_X�g�h5uhy5�~C�If�4G�<ƖPR�H� $N>-N8HNCKN>_N@0R:TC'T@�T<�TC�TKJU8*YF�[<\>1\: _>U_KdK�e>�fK	g:@g<LhKfk<�kF�k9BlF8n@�s1�v&awF^y@}�Kp�C��@̑:�