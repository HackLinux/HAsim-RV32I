G~5L0D~0E�3D}/Es'7U';g/F-B.Fv,Ef)<[+?a0Hh,Ad.Ah3Jo4Gn0Eh*Cl(Fh'B]&>X'<_+Ee)?c(>`%8U$5L&8R+=W.@X5Lc3K],?X2I\.CT'<K+<Q0DX3CO/;C'5?*5>*3*117#6E&:N!5I*;'8(< /@+>O*;D)<G&4B!.=#09!/; .<!,=-A/@#5E&6J(8L%7I#5G86>:5$B&?&B!@:1,,2 0*.2+/231!7!)=1/#//!0!0$0!.#;!+C#-E%0C$.D+5*4)5)6�-=+?*?(:%3#.!#9! 6!0  2."-D*9P21=S.'?�",B	8,- 611"5 '< 97� � 2=>4>@4?@3@A6CD:GH:HH<IJ�>IJ>JJBNLFRQESSFTTEUUEQUETUHWXIZ[K^_N_`OaeM_cQcgTef\ln]mq\mp\kl]kk_onasraurasq]no\ln\mn]oq_qs`rt^rt� � � � � � 8FT9GU6CR5BQ8DT6BR8DV9GY8EV6FV7EU4@P6BP4AP2>L0;H.:F/9E/:C-8C.7@+6?*6>)4;&.6"*4#+3"*2")2$,6"*2�!*1#&-BEDCDEFHHIKLKK2: ;75#<:#+G (D90#'A >"'B(3P#-M"D)E+"<7�";{!#;%,A'-C&0D&+@! 64 "6*3!7"8 !:%-E)3I!&;,7P1<S07 1<!3=!09)-,5%29!,1&0*:2C/@+=+;29-*&,(1,0)/!/5 /6 /:,7*0-7!2?"2>$5@2?%6C&5>(38$-0(+(/80=,;&2%0$+" $&) -4'8A#8E 3D!3=34 04,2*1"0< /:!.;!1?#4=!2=!/=!1? 0< -:#/;$0:",2!.5!3;&7B&8@#7G%7C&4:%5A!7I":L%;I*?J-BG(=>&8:*46 (,"'''")"/<'9K*=N);G)7?'27!01 22"-4.</B$9D6<+4"2B!4E&9H"2>$8B�"5F
2?,2+4"2B#6E!3?"0>%8I%5C(8H(=L�&;L':I$6F&:J':K"/>'5A);E!5=/7%6A!5E':G$5D*8@'6?+>I":D 6:"04$3:%;A%9A+=I);G+=G/@I%1; .<#5A'>Q&9@'7=&:B/<(?P)=I,=H+?G(6>&/6'/5%/!-;%:I&>J(=L*>D57 .2'-#(,5$9F*?P'@S(@R(>P!5G+=M*<N*?P):I):K(=J'9K%7I&9J'7G&7D(9H'<C'>?'79)6?%4E"3D(;L,E.>V+7Q'2I2?Z0@X+;Q(5F"4:$4:';?$48'6A)>K"5D#:G&@L#;K%>E&;B"8B!5;3="8D%:E$8@$7B&:H$;D&;>$46%27$5:&8B'<G&9D(;L&9H*?J(=J%7I':K(:L&:N#8M%4I#5A%9?-3"2>$4D&3D"3B!1?,5 /:"/>&4B&6@ /:,7-;+6*8 -< /: ,2((2=B1>C0>@=OS;NS<NV>RX�?RYu?S[?SY8EJ:JN<LP&?#)A%5;&9>$5:$28,5*7$/(4!/=(;H';G(@F04%15'39$9D$<F'<M)?O'>M+AO,@H%37%,(1-6+6 1@"8H$8J$9N&=T)?U-DW0F\/FS+BE'9?!59 -4(7@(7B);G':G0ET/CW-DY-FW#07!+1!,3%4E0?T8J`5D]?Sk7Mc/F]*DX"5H+? 3#4$2D$6F-;5>(5-7+4,5'1-7"2 ,D*9P'4MGp�R��Y�C_wC`w@]tC_u;Zo7O_2AL$4B#19#3=$4B&8B&4@*;H';G(<L*@N%8I"1D'6C!1C!2C%5C#4C$5BH]dH_fF]dF^dF_fJaj�JcjKbiH`fF[`F\`�H]bG^cDX`F]f$4F&9J'>G:<#6A+>O/DO2GR,BN(?P1IU/IY0K\1JW/GS->K-;C&9>#3;!3C(?P.IT&AJ-IO3JY2I\1IW1K[+DY/Ha-FW/F]2Jh2Nn3Oq,Db(:T!1S(?h-Ba-7M.@d'<_+@u2I�1H{0Dv.=l,>b+7]&4^,?v2H�5M�1E�3F�3I{4H|4G�/C�3I�-B}+<y/A�0C�):s+=o0Ev,A~/F�-Ao(?h+?]1Eg1Hk/Ga'7U4Jx3Lq,Gl/Gk/Fi)C]'=S%8S&@X&C\$:X#:W$:L#3E*=Z.DX&6J5La,BX2I\0EX*BT+AW.BX4FX2?H%/;)5 *6#/&1*5*=P&;R%2K"2H%8I .D#5G+=G)7=$3<!-;"/>$4@"3>!1?#0AY*:N(=L#7M'8M%5I"3F$7J';M7;@:6(E'@$>:1/--3 2-230/!7"50"7 '</,$,/ ."0 0%<!)=$,B%0C%-C+3/7*4%/,4+5,:*?&:#5#/!3 !6/'%3-+-5M$>#-E%3I *@ :!61!<"=#:!*=,6F-6G#-A:L^0@V-;M1@Q0>R +D(B; :� � 2=>4?@4@@5BC6BD7EG:GH<IJ�@KL>JJ@LLBOPESS�FTTFSTFUVHXXJ[\N_`QbcRbdPbfRfhVhj\mn]oq_qs]no]mm_ooasrbrrasr^np�\ln\np_qs_su`st� � � � � � ;HU;IW:GV7DU6CR5BS5AS7DU8FV7GU7EU6CR6BP4@N1=K0;H.:F-9E.9D/8C/8A.8@,6>)4='19$,6#+3")4!)3"*2�"+2"*2")0DECDEFHJLKMPQN0 :%=#=!>!9%A"'D%-I$C4,-3#(E%.M'H ,N/"8021 5#$9#$;#'9$$8!57"#<36!4!'?"%>%*? !:. %<+0G 0:!1="6>"3: 1:!2;#4; 16,9/@-C/A.?-<)1(,!)%2,9+8 /:#3=%4?+4-2#5=!09"2</CK(<F(9@&28*/)+!%")-808,2&,$+&+&#!0;%6C#5= 2>,7)1(,$& $%,#3=&5@#3A$2B"2>%4?#/;$1B/=+8!-3 *,)*&( 04$6<"6>/"7H%6?",./= 8N!8M(=H(AH*AD"21$0/".-++*)#)*4%6A'8G*;J(:B(44(02!,1 43(/*9"5F%8E!39!0;%7E%;I#8C!3=#5A!4E#6A01'/"2B"5F"5D%8C%9E&8B-BK-BO(=J�&9J'8G#3C$8J&:J(7H-?C%4; .2 *0%6A"3B*<H(:B#17"28"3<2844 .6 0<"8B!5='7C*=H*>F'9C(8#3C$9L#7G&8B(8B%6?!2=&<L&>J,?L-?C&24)35(04$- 1<%9C(:H);I(;B 46!/1).-5%8I*=P*?P*@T'>S$<J 4: 6D):I*=J)7?"4:"6>"5F%7C"2D%8E&6B+9G0GL)>?)9A ,<"3H&9J$9,<R%/K"(<%-E,9R)7K&0@,8L)3O(.H,4L1>U2@V0>T#,E 91*#$3#)=$>#>#?#? @(G!/M&6T+;Y1?[0=X/9U+6Q'2K#,E!&?84" 4&(8(.>'.A'/C'0C&/B&,@%+?&/B+9O+8Q&3L"/H+G�%=!-I%5S+<Y+;Y+;W*7R'3M",D!'="7#*='0C1=C0>B0<@=MQ;LQ;MS<QV?TY�>RXv>RZ?S[8FJ9IM<LP*6N+9S(0L$6:$16!+1'.%0'0 .:"3B%9C!3; 12/2-52<)=G(=H%8I%:I$:F(:F&:B27'-&2/>,>/A3B4F#7K&<N(;L,CV,DZ(@P%9?!15,3(2#0;(:J+AS!1=+>O2K\,BX"-4%0;!-5%0;.@T4F\1BW*=P5JaAXo/@]%7S+;%2&7*=N3H_3I_1?W1<S&2B%1'0 +64ER6CR&2B%5$<$A!5M6Vn8Rj;ZoFc|A\u9Pc7Sc/DO0?H-=G'3=*<F'<I"2:*>F%7E(:J*<P&>L#6G"3D#3G 2D!3C&8H%6E&4BEYaF[dG^eH_fHahKdkLfl�LelKdkH`fG^c�H_dEH_b?S[CW_%5?$1B*<F'8G(:L+AO5NW5KW0GR+EO+GW)F])H]4MX2GP+;C%17'. .:$8D/HS'GK 2<*?J4PX2O\0HV+=I*@R-E[1Ja1Ig1Hg1Hk2Jj/Eg2Fj,@n-Fy(9`,@d):Y->m,Av0Ez1H{-By.@r+?e*9d+=o4H�4G�.A�0G�0F�1O�)Cs0G�0D�3J�-A�0B�/A�2E�1G�0E��0F�1K�.Ar#7_0Dr-Em2Kt+?c-Bm5Iw3Jq0Kp1Ko0Ij-Fe%?W"<R)DU%>K"@P1B".B/D_0Ib(:L%2C*=T-B[0H^.AX*AX+A]/C_5I[1>G")4!03 )6!000E%6M%:S)>U*@X&9L -@$6D+=E+8=%/7'3-=$9J7> /:%2C(9L'<M"4H%6K$2F%5I&7J'=I'>A9=@;9(A#;4103433 3- 3 632)=0/2/.,(00#0$4#8 &:!(;#,=$,B-7-9)5$-*4*5*7+>(;%6&3#8$;5!!1".)!'?5&*.$+@!5!#?,7L4@T5@Q1=M*1D '6'5K#3M .D&4L0>R/>S(F&A:"9 %:":'/?&0B!5%6(� �  1?>�4@@5BC6BD7DE:GH;IK?LM?NO?LM>MNAOODRRFTTFVUFUVFTTHXXL]^QccRffRefUgiUgkXjl\op\pr`tv`qr^nn^op�aqqasr_no]mm\ln\mn_rsbvvatu� � � � � � <IV>KZ;HW8EV7DU5BS4AR3@Q8GV�7FU9FU6CP4@N1<I0<J/;I.:F/:E.9D/8C/9A.9@+5=)3;%.7$,6"*4!(3 (0"+2#+1"+2#*1FDDDFIJLMOP STR")3$9%A75. :;&&9#/Q)7["0R1-0(#  6 #<80 9!$="%> ": &>1("&<#%=!!5 $<!%=33/7 1: 26+/"3<#4=%37.5,>+<.>1B 4@/;-8&1%1(7 /<!-; -:&6>'9A!5=#4="04%-#2;+=E)6=&26#,/%&%%#%!(/8 4:!-1&+%)*+"' .6 2>$5@"-4!-1,3+1>&+"(%+)/"0<!/?%5C!1?/= 0<0?/; /:"/8#-/ ((*()),3(:B#6G!4I#8=%).>3H'=K'<G';A%9A%67&34$,.+++,&-&8B*<F)=I*@N,>B)23$02+2*.+2 1@#5K#8K 3@#4C%6E"8F!7="2<"6F2E%2?"08!-;-:!0=$7B�);E*9@/AK*>N�#6GY&9J):G%6K%8I&<H'9C*8@%17!,3+;C0BL)<I':A%59,0"12,228/42?!2E"5D&7D.BJ,@H)<G%6E$5D$;D 5@"6H&;L"4F#8G#8E"<B'>I+>E%<?%96'33()+1'8A+;C*8@&8D'9A#39)7;,4&6B3KY)>Q+>O'<M%;I 5:*1#7C':K':G'29(6>*<F0A 0:*9D(:F)=G:MT8NV+=G"2>!0C&9H *@�����������������������µ����������ż�ʁ����������������
�����������������������³�������Á�����Ÿ�Ĵ������������������������������³��������������o��OhoD\bDZ`CW_�DX`�DY^CW]@TZ@T\BX`�D[bDZbD\f�F]f EZa�DX`�EY_|EZ_DY^CY]AV[AY_DZ`E^eF^dD[bDZb(*"(.&3*7"2>/7!15#/3(.*4!3=)=I(8F$4B 0<!3=);E'8A!29-9/<0@+9)6*;/A!3E%7I'9K(@R)>Q&9H#0=$.:&3>$4D%6E&<J(;L%5C*?P1H[-DW".<%1E*7#/C):S0AV.AT3H[.?T1A_%0S)J:*=&5N7Ka7Oe;Ni2C^/:S(0P'8".!)5<JZ=K[/;I!1?'9!=$@,B;Uo9Tm?_uDYt9Tg9Yi.@L-;C,<D-;C%:?/8$7B(>L*@N(=L(;J$7D"4D#5E"3B!5C 0@"4F#2C"5BE_gF`hG`gHahJcjKemPipLfnKemLflIbgG_e�H`fI`eE]gD\f%6?&5B�):I)<K(=H3GO4IT/GS.GT+F[+Ha*CZ6KR)9?"48".2!)%9E0HR0LR*DH%9C.ET1M[*HR'=K$5F-BU0H`1Ig0Kf1Ig1Kk1Ge0Gj1Fq,Bp(<p)>o/Bs0Dp0D~-B}0Cr,<n,<x+@u+?m+>m;T�8K�6J�4K�/F�0F�/F�*A|0E�/F�0F�%8u,@�0E�=T�9M�4J�.D�+>u0Bt-Bs*?p0Fr1Jy4K�0Ev1H{0Fr,Dl1Hq6Qv/Gg*A^;I'@S&9J!8G1B 1F+?]2Jj0F^(=L':K.C^/D_,@X(>V,Eb1Jg.Fb3DS.8D$3<",4(1(4-?%:O(;V'>[&>X*@\&8N)9Q+>O(9B%/7"/8$0:%4E4>36 0<&7H*=P#5M"4L&7J&8J+>Q-@O+<E,<B�:^="B: =&>4167::!;421#6!7"7!8&<+/,+//,