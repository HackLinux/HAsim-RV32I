t[�U���    t3�t�M���   �������
ǅ��������E���������   j h�   j j ha  h����UR�FU�����E���   �u  h(  j ������Q�"o����h(  j ������R�o�����E���   �Q8Rh��T h��T ������P�MQ�"����������������� t�������  �U���   �H8Q�UR������P�MQ�4����������������� t��������   �UR������P�MQ������������������� t�������   �UR�EP�I@���������������� t�������o�M���   �B8P�MQ������R�EP�N����������������� t�������4�MQ������R�EP�0����������������� t��������������M�3��Sk����]���U����} u
�z�����  �} uf�} tR�E���    t3�t�U���   �E���E�����M�U����   j h�   j j h�   h����EP�?S�����M���   �o  �} uf�} tR�U���    t3�t�M���   �U���E�����E�M����   j h�   j j h�   h����UR��R�����E���   �  �} uf�} tR�M���    t3�t�E���   �M���E�����U�E􉂀   j h�   j j h�   h����MQ�gR�����U���   �  �} uf�} tR�E���    t3�t�U���   �E���E�����M�U����   j h�   j j h�   h����EP��Q�����M���   �+  �} uf�} tR�U���    t3�t�M���   �U���E�����E�M쉈�   j h�   j j h�   h����UR�Q�����E���   �   h8  j �MQ�nk�����}(}ju�UR�EP�vA�����h  �MQ�UR�_A����j�EP�M��Q�Z����h  �UR�E��3P�Z����h  �MQ�U��4  R�wZ����h  �EP�M��5  Q�\Z�����U�E ��6  �M�U$��7  3���]������������U���4�E�    �} u
�z����  �} uf�} tR�E���    t3�t�U���   �E���E�����M�UЉ��   j h�   j j h�   h����EP�8P�����M���   �&  �} uf�} tR�U���    t3�t�M���   �U���E�����E�M̉��   j h�   j j h�   h����UR��O�����E���   �  j �MQ�UR�l;�����E��}� t�E��  �}}e�E�    �EP蒋�����E��M�Q�U�R�EP�MQ�;�����E��}� u)�U�Rj �E�P�Li�����MQ�U�R�EP�H  ���E��)  �MQ�UR�EP�D�����E�}� t�E��  j�M��Q�UR�EP�B�����E�}� t�E���   h   �M��3Q�UR�EP�uB�����E�}� t�E��   h   �M��4  Q�UR�EP�EB�����E��}� t�E��   h   �M��5  Q�UR�EP�B�����E܃}� t�E��S�M��6  R�EP�MQ��?�����E؃}� t�E��+�U��7  P�MQ�UR��?�����Eԃ}� t�E���E���]��������������U����E�    �} u
�z����c  �} uc�} tO�E���    t3�t�U���   �E���E�����M�U����   j h�   j j j;h����EP�{M�����M���   ��   �} uc�} tO�U���    t3�t�M���   �U���E�����E�M􉈀   j h�   j j j<h����UR�M�����E���   �   �M�U��j�M��Q�U��R�bV����j�E��3P�M��!Q�JV����j!�U��4  R�E��6P�/V����j!�M��5  Q�