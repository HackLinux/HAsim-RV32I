Ji?��X{�����"k�N!�|,!jE�G}���T��"a��=��W1�b64�_�<ZYz�-�9"x5=4W��U^R2e�T=�j�:��w��Ј�����ۺ�sOSc���TOE�1��!�"���V��;?�)��n�O6&~�OK��u��_�C���ߙ>�`L�&z��C0@⸧��,���2�4��r�M�F�D��g���:�wJ�S�5Z-�_ά�!���宙��LG�G�v:ײ��tfs��mg-	
.M��Ф���F��s�.V}�T�]y�w��_�
��j|9��ըNaB�N�7��d�y����G�kgC���K�nh��Ì�S�i0� �]俅w���Բ��*<g���ɠ9%|YRA�9?����r1aӤջ��[�Pq1-��枊I��$ �Q�aֺr_:L4��k"�dh�/�v��R#���<�l<��h��KN��|s��ꚥSb��ũ_�{L[�䶩�����gM��H� �dv�8t��v�n$�<�� ��2��Ғ�$�;'6��1�1�o�f�MT�xb��m�?��Sw�3�@3���BO�����_/��_5�8{�G3j�kn�PkIĖ{\�A��L�P��.B�Zv��%RE?�XCؐ���	�	j��ƛ�W,���������j͋x�N�W�I�s����; ��@����������.�t��}�K�K�E~��H���<�=�N �D'X��>�%���̣&��|k=��Bh��9Ϲ�F�<v�Ғ���&��a��
u�ܮU�}����
��35
�zk�{vvw*�j�Q6����&����r����ћ�c�Gy�g������~G �l��8�(4�P����H���)��o��G�Ĥ�A��E X
G*�r�-_�iڔ�9S$V�� r���
��߯X�j���Yd`�z�B.�KV#���t��j�!�%U#�f�ʽs:�E���q�D�&P���	�NL�O<�/�1S�Vɽ�e���X����J��n�����'��fS�^��V�a��
��P���|{���bS7N@���㠛;2�F9 �3�6���:
�7�����χIo+�,h�
�!8c�B��	�	|Q���ˇ�C.�I7�U�F�ϛ���X8ƿ�+xt��������	j@�l'�!)0)�V�C��+�_��dԠ�d�#������H�OR٩p��5�{V�̲���O���뙽R$f�S��(�ƂSmSߺc�I�����9l��l�@q;�H9��r��.���!��B��gv*�@�,D��aٹ0[�l�΅<�Y��&<��ҵ���-=K��I���]B�|�����cE�0�tT����{�!��+�qI�X�9�|$.x+�Ţ�E�O5:[���S�0��u!�j[|�Le5҄+��0n�ߓ�?v"��ųc�"�52��x�w(	�$}i�»�������nю���X.�ҳk:��d���)��zN�=��^�\A��HG������k��]�6	6���̎����V�J}�q�^�_�P9 �|O����<���������:�i��*��r,���Bx�̛�=9<���1X�������Y�Gʑ���QC55)�vB��Rߖ^���гK�;�a��eHNQ�9	�?����d	�tD]V|1���. ߒ�s�lz����fz*p���v���$w�3�2�e0��E��C
���<�h�p�"�G/;��sb2�(n	U��t�����ٞ�Ϡ@EI�Hlh੨��m 1:g^��qU�g`��J�X�������:�����9��=C9�K`�w�t�h�[~��c�7lC��ZIbTaf��g�
�n����(4���Љ��Њ�w�s�	W��韵�N��0|�>0��? �_�7Β��lZ+��⑜�3AZ�����#_m����������e}$��꼂Ym���K�@|E�
ְ���7�˅�i�IN�XB���*�u�k�X����i`Xw߸�!���7e��_�&�h�����'bhV��г�K���k��|����1��	<X��<d��uUHCHbQீ4kp-�%��2r�#��4�0�|E=B�Y�
s��Y�|��W>ߺ�w)�UU���V8N��leN��o9-A���;�A��@ܶ�琂NI�U��}1<~+�8�q�d�Y5R��-u���_��1�D�w�y;����l)��kJ�F��a-�d�����tl�~r�g��]0I4�$��,���P�1aP;���Qt�R�蹢C%`��q�¢��:,���G-���}0��9��d�m}ݰ�-�e��ޢR)��د�s���%���9eJ�ym�!��*���[�C�:����J����>b��8+{.ӒvJ;u �m���Ew�&��S�+�*=�O6����Y��>i�g���n�������?�'(�l��v[�XF�v���2g�<4���c����k��ڋ[�������;>ip��0y�G������nd��i[W�·L~�	�5|��Ԩ����8	�H�U��հ}g����}����۝��U���ј�����M@z�S��F�L����bd��~��G��-�*�Q�T�2FY�����0:��6������%;k�l'��\j"׭�@�[����Q����G���q����(��9�B{�Ht(�ߒy�1Ε����?v{��8�����<]@��Z$V1��h���芙f�D[��]ї��z��#�g��i��/�z&�6q@?�X��Eg��0R�꾰-��Vu�K����|F��~����t�v�hIJ�����#�f���ކ�V�%������?�#��dzZ�<	�\���F�6���ઓ�zy�?�΂e�OcC�|���$��)�9���Z�z��p-�	[p#:b]4n�{�O�YȘ�����W����Ȅ�$���+�����)Q.׮�8/��ה ,���T�������"M���4Z�P���h�0�g�,�(_%
p�;x�s}�GhE~r_V����!I��L�r�~����+�J޻zD��cJ�<�3�qh�Ib�6�<�ʁ$�?�ձ����܊8���l %�G
.$�i��m����[����h6Z]���c�tQ�:a}m���G��Lˌ��u!h�7��*���+�Y����|h��&��f�L����m[ԋV��)p-#{��О�ܯD�h��.{�-}]��0����?��$^CWa��y%xo�݂�k���?K��<��i��I��)�H,��]q|	�/�]0���/�i&6�
w[���Z7�.TJ���㾵��JF���ܢv�#��z\w�,��F󻊎�e��B
A\��M�Tĝݤ�\��1�Ő�hp̏P�[�D�,���+�a�S�5�t*�~0`�^���|]\g;͐D�sM��"�kwav�h�V"��J_��9�?/����!_(h���b�����=cL��衳��R�Zg����9�Z�8B`y{���Ÿ�/%b������z�BYw^G��ɤ��8�Ӂ�����-����'J����`�sZE���%��iŇ������^&�9�A����W�cl��=�]��������Mj�t$��ZD[��(f~�qMNK�-g�
��?:z\F7Np��ˈ�S#�?z}�&؉���E��Ź�	��Il�(��0>y@�|_��f���g:R?=I��a+뭞<�����ܸ���|�+��6>PvW��6z�J�me�2�z�O@��� i!���d��T�HK��.�N�˔Y��O�{�vB��C���*�Kfd�UZ�4iT�2���B/����,�;)�_� ��
?����w8��)
��9;I؂��'�DTx��M�g�?�n$F�\��
����ol}Y���_��of{D�,x��������h�/��Xе�=}��;�QP����l�A���i�zS���G�Z�
-?��:�Q�'�f�;;��.(t��)��j�v]x}b9�F|�x�@�z�RE�d�t��~�iZn߬U>+�1s2�4�|$��Pm�z��Vu�����B�;��%�����g�}!IP ���u�?D�A���M�%(=�`1�<b�ؕ�t��ǥ������IOW2=�Sm59�q��D�,ReuT94;��m~L�i��u�r#al�������ze?�u�>�C���m�=\�=�<�]��g�^��wvBz�FT�e5�fu5!��
��'S�nFh'EWǥd��S�C薪fl'w��WTW:�������Dv�7�SR{&��*ߌ�{\�-��e�X�Y�gcn�J��;,'}�k���(�6�R��<���W��Sw����J@������I�|��s�<W�U�42�Ir����^e�b����$��+O?�|S��L��Y�H=�z\�:�QUԘDÓ�@A�V�
�����؇�L���T�!sr?��4�^���>a�������7�d,���E��}�+#u e�tʦ�����ݭփ����Kyt���+��7gSh��v�~��W\~�U��iw��p~�y�������"9z�j,\��'�{��H��r�l����@Ҙ6V��q`S|q�ȺSS��1>��Q�S1������z�6Ƨ�T�U?�9&_�X��t��V�;����ņ{K�I�F���Yt�A$C�\�;"�^�������'��jѰ�_H���@E뙿�����s��Ԝ��n[e��YD.V�d;�on��b����1��
fѦ��+*��R�$l���fx�r@㾞{�x!���d��R�y~0��Jk~f1�,��+j�42ƍ'%}�������z�<�	o�J\A˔\�Eo��|��Z�s�X��&��zHa!1���	��U{A䧝w**��]�2�i����U��'5��,��\8�Z�}���;�NV_���#4~�¦�����L�j��7���GY�Ƹ��o�.-BĲ�5yɥJ��/�\?)�GԷ�bA��w��?�^bJ����h� �����r��5���@p#`8���3uE0ui�|�q�Ω�ONd}�Ev׷��:?m��F/�B�6o��[lֺ�ԳN�/��ǎ�7�|WFS=u���k����$�N*�/Ԙdb���D\���\
�Pl�ێ��Q3�2A}`'!��J�m�`"�{�3�zg��#�	�eS ����r�S?���/��]����Yz�Z�oh'�.�4t7�\)������+ 嵽��.<>���F�Ć�e
��u$2�K��A��g�� yԿ�HS߾e9T�Nyʯ����DG�ÉloQ�Hj�5}%�
<S��m��%�2u-XH2�ӟS����O��Ls��v���N���/�J�~tߣ~c����i�j+����$�}6���ы�Q�H[%�l�ۅST���0�H���H�US�F����ys��8c_	�ǁ�x7�O�/����P����(�l�}�'I/<�9�%!���h�/����P�L����C���W��ۊt:*��
�zb���h5����r�҉� |b	fD{�u:�w/xDN���0s����0�L�+ar��u�-�1y>Q着�}�"��E�o=��~#g@]D�p����Q�U�9�N�����+�ޖ�ٍ(�"��t����	��
�h���*ũ��r�u�V�A�3O�Z+`��%`ff�#]f���w<�o,�7.I|�\��up��&���% p�0�s�2�ڵlD;sC� |���+s�ʛ�Y�N����lr�S���dl!b5�|����i�k�K��|z��P�_�zOpV@�(Z�����l%p��-��LIFM�4xnQ�j7�\U���3s�/b�p�P-���a��_rƚ� `�4��VՖt���� A�Ny�pZ���MkQ�娅���3zl�ޝ^xכ��?:��՜J�9ݔ���x\�>W",d�����
Y�,��wƶm
h���%��3�r���-�~�DPaJ}����	eiǎ4d���`>b'��)}5!�c�h��C��w/���m��� 8�P�d�#��y����q[�;�f����w�A�	����>�#7H���?-���r1.؏{���'��s�%瀺p��T����ܭb�2��Z�Ө�+����ڿJH�3o j�H�.R��ֱ��¶��ɝ�u����.�RƌG���P�V�:A<r��o5N=�}���(��f4�j}����~����g�Q��b��7�#S�eQ%��|e�HR�s�Ͷ�X�._�{�M���#�@ KY�a���_�i��M��q�]_�^���5�U;���#�y�x�.H��~��%��+�P8b�j��
s���h	�Ffc�o3V��n�ȹ#�Fn@]�gP�}�4����[4����
W(=�Z���W�cȫ7w�D���l�2ܾ��WLٯÂ�I�~<Sr��U`��BOB�%Tu�9���&w�$Ha�K���p������W�hxڈ��S��w!�`��l[�Ϥ��(te/�	��nLq��z�Tɢ[��ʉ��χ��+8*���%q�ONu�[�w��!�4ŏѶF�L�'��A���ؒ?B�H�qy�lv	��?X�T�����HT`�%�I�VC{C��P���Y�;%��V����]��2���U~��nϘ��H���`���i�g�
XQĈ{7���s���E��d���qva���� �u�r,���l��#�KX ����'��}��t�uI��'j�	A�T�����}F�x��җ�.�,K�r��
�(5���!i���d���&%�1Owb��`&����Ψ��{��XBeĻ�ʐ��!���65J�#r�ǟ2Q
6�*B��w���䚪6��˞ot��찝H�Q�:>�^���I����S)�i���u�ak�=�DzV��=ܢ_!f��]�����W�sq����^^؇�����!�>_U�3[9`^��SC�2���-U؊hl�g`�MM����;Yw�{�ǹ��*��(��+"�k-G�&���)�����e@���}���"�:�<?�.-ٱ)<D���^&�M�pPU�� �
�z�]0���1��;��0�m#�q�q��e����F�s�('*T\�M�y���N�vN6)[ƹ��/�t�}����.�����;R云I�Lݑ�-�����(p����N�Jn�&tT�T����2T��Q�I�I��39��#*�Ȟ�n,��U�W��)��纤{Q�O�l�����9v�]���.H��#p�= 5�v{���}��l�Z���df���������r}�4��޸3_{坾 f�|��2�{ޞ'�<���zp��8WT"�? ͉p���O7M���7��`�+��\)%��䆐���J�ٚ���$k,�f�����Z�W�0�9D[.��8UP���G���S��5�8|:��J��hT ����|O�Ɯ�{��L,����$2E"�*����ЍD�W����u����ց�/ٷ�%6����+�L�5�ްT$�-�.�%��{^���'���^��]`���p��G�X��X�����#��^�,=0�%�B��i9��%b�\(�pc
꾝ߠen��Bu]���_�dJ3,ܗ �Q�8�����������'��GQ&R��	��}�q��Gi�����7?��"�Z~��\�adef�ԛ��K�_�Nw����:,�����]#�i*�Р'C�r�A�~4����l�|]�7ۃk�s$���hv��L1x˅�1�V�,j��

��Q��2�Q����u��%�;��_��G�\�yʏ=n���';V�Q[έu<�tK+��~hX�&{ME|;7���݂pˠQ�Ju&�w��D%/ԭ�դl�h�^�m �35���ۮ�'d���y}��XX���??|^2����������ZG"���l�DC���̽n�k)�5Zm�+��Nױ8S�����r�#���(Bٽ�.k��Jy#�7~hz�Y^Kn�.T#i�K�
�B\� Z4�F��ęl<�ٛ�y����4ZM+�gW�Αh�4�j�Mץ�$~{r~�7C�n�!��4��
��ĳ��~�����&%�RL}/�m'�R�֏�9B���&����ʍ�m�����-	�8�4��������(���q+71��V�OT�9U7�R�찠na�JZ�5���zl���������!ݏ�TĮT	�	�l��p]��WK����I{����[4�Hf=��vk<����=��J��4��S���=���yp���O
���A��fO����l����+R��L5vL���a�[ʰ�J	��m�l��cb�,���n(���ҩ����K�&RЭ�3\�vcx�a恈9�AɦX~ᣬ+����$Ɋx�H�}#T_����lϿ�\s�/�3z�)�_�Ǣ]�>y�	� g��I�5��ݠ�3� �_�����CX6�D��%7�����2[����F�}��Ɩ��m�~U\��af�Wv���?���آ[�:p?ٖj���Z�k��I�����<98|����I�
��|��W~����}[�������~9��t���y�S]ݕqT�1�[�u�Fj(N�=���#�=��l�����S�:�Z�V\jL���`�W2���2ij/��=زr7��Mԡ����_�M���FX$E��H�5S	���OD���K��T|Ў�j"R�K�1y�]�����!Gu ���El__���9�'%�����CQ���'W��Xx��ϥ��w�&A����͌�ʠ�ciIH��ױd؊���!&ǩ�Y�y�$�L�Qf����������en���m�=^3J�k���A8}���Q��;��[���{�hDw�����+�еO�xnO�-XS"��>}F�SJ��]ў}݈��]Y�TX@�*���Ɂ��J�'��^11�\�L�RJ��j��U�dD�]���3�c��+BC�f�V*�����4����@qy�g7D�w[�}���"ԗb��n��
|a��	�ӟ]\-m�#���/T�i�>ad�%��_cR��B�H�);r���ܣ��'�\���3��q�<k�ڭ�C�X��#�O`��4�Ҋɻ���/���,!/S��
׋l���=K�dU�jn��,9�>�����8�+����.lg�ښ��Uw��.�X����x���_B��He�M�y��c��d��D���0o9z�o�b����ƔWq���~���}�Jަ���� e���n��������P�ʴ E�({ྰ����k����
�����É�o��"UUk�I���:Jfʝ �N�Jv�}��:Vĵ�������X�I��q�\T��4�&3Q<�__;���텹��Fl��~[��F�X�Jp�"�$yd��zX��aB����p�]�@�Ȍ��*�0�v�5�w#*��脇�rt!��K���]��{�;�"��B8���L�<��"��p�Q��4I�U;�)I��>�'���z�m�?DC㮷�zBͿ7��Ѫ8��I«��e�x�}� �{�Lv<�chZI6��ȏ��V�]u�b�N�z�C�r�3�̣�3a�jNd�B�>�뤻egB}+�n4`zj�\�g�=D<�����!~���Ɨ�c%��R�z�t��udUو�}Y��Jl��	ٕt`Uls�Tqn�'��a�=�[v����v�*�#�=�蜂ċtW:�kl�Ħl�b2��됞Ў�%5x��2����
�@����q�x���a��~�-,�;�� a�"�&l/��C��>�%���l�=��'&��?iJp�+�c�$�R���7�v�	����2���}�����4$ 'iqd�b�e$2�����cJ�@�h��bp����6����U)�v�/�m�WsP1M�o��/X�������K9ʹ_La�0���$Y�B����G��-�HL�y6��fx�zg��ɋ�l#@�E��J�nG���K���lcL�{�k#��FX�M�čx����t� �����s s�a��CK���ٰ.�b�hz	}Z�0�������&���׃Ȑ��zS������8��r#5̉s�#_�Dە��1�2>e���_.!��^Ѥ�71��q���R���(k��� �zj9�t4eګD%���Q�ynf�z���,�� e���[:���;8Ns�_d��9�U�2�{�g���>O������� ו�у��N-���Lp�
dw��ϭ����=�^;�n�m �i�r�銰���o�	���c]�O�d��a��3ܝ���#�X��]'����o��h�vo:p&ڜ�$?~'{�~�ZV�{k��'Wl��%d��ӍRY�H��[:���N**��PG�Hb�F����p�G��/5�%���A��bw6?g����w�6���&�����yԶ��	g_F�8���8�CO��<�����ܭ����f_�Ve+q2U�O�OI�~���T+q|u��S�F�E�����k�"@��SX�`�F����+ΞʇO��߅-�[��'\��Z�p��G���J&KG[ ��=��D����!�����̦n�'��%�P��W��k�<�4�6�c�@�'`{�#���	0�(�Z]_c��
guz��y�-�ˍ�	mfq���/kXw��!���)bܷ*���࿇��n��H>��ogNN2Dk�����o�}�]��߄��G��r��u"ӕX���8A���(NU���H�`|�KN$�oAƅs��1���­�I����C�n�����Z9���d|�9�<����묂o#&�oɱ������/𺑬����K3Ĝ��uW۾<3�?�����]t�8ZP��I+9��W�!��+�q�e $r��+��y{E��*B|l���r�x���g�rV�&;�}�Uf�H��dj������|S�M��[��32S�GD��Y����x7����mۏ���!�y����g�S�0�D�Q)�(�� �4���N���(�Υ��Z�׬C�=Le����A|,: *Ʈ$,�g��*��7tY�se�T�]����9��� a��^��	�Zб��J���*�鑽q��|}e�4�	:�7�� �9j+��|����c�%�7h�