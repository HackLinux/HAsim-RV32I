�`��P�W�f�єl�n~�� ��U�S��y�4���
-(���//`�O�4	<̌�3]\1�u���Z�:�ㅜ3�V΁;ST�s��L��j=i��A<�n4c�/p%�L\�[�v@�M&� 7 �]@���@A�n�?/Y!)��{н;$��1�>���Va�3�M���7:��9,�1=0��`K����0���qR;��Q�'�P�TGP)ǀl.�)����q�g�Q^��v�J�-K�@�AA�МX��b0(���O�t^���A0��;\pq'�bN��;�%}��v7I�\�e��
x���K� �j7 �K��  Y�����Ԍ�
,�(� ���]��� 6+�y���wA�txo���\����pj[��
�\1`���vϼO��]���( �0�v��6Th�i`8����� +1�� � ���r
�&Z��&A9���. jA��O�}߽��_M��Bs�,����]��S���ݠ1�O��� �AA�ͤvB���Ā�� �(���
�� �� ���o��-�1#X�/,��0׏4N��N�<��+��`��P5�2�i�3"�
�
B
�Bl�!��R  ��6�� ҩ�p��� �� ��b�W0]p����9����ȹ0D�ꋠ�M������h$ ��"
"
b
�
��L� �  A�� �o�&�� V@ �$ ����� �
�BШ �� �$ ����Q1Uo#MrJ�v׮�����p����x�,����b�	�a"�
"
�
a� 
�� )l.�v!�	� �ą��BB�	"P� �� ����������i���.�n�ΪJ���1� ���  ���
Q� ����� �2 �./�
���o�@ �
���T
�B ����� �a&2e&k�O������AS�W&��������!@�	�P��#b��� �� �H 	 �8 �+Z��G(r�,��-*Q&�=�S�x�.�/�(2�.��(�$ �38��
�2A$���131s��د�'�N�FN�J�i $�s8�R�1�A43E4sI4�L:.��U�n�?O7����2N�8s=�O7sy7�}7�8"53VN�]-��\Sh,�4J�o73�:3�:s�:�����XJs�2R�'s19�m3�U7S�<��=3�=s���;d�;�A�c.���Js�<��?��?�@4 �&KSU;S�C�_3)f��jM��(�@t-B�1C45Cg�=�t>��6D�2�"L�'S?C�YE�]E�aF%�C��>SaDs�D��E2�B�eG�H4�Ht��t
8T>�F�N�*N�M<T%<�)H��J��K4�KbkF��I�EA�HN��?�7�K��Mt�M��H4�L��'3�<tK�y ��Ot�O��O�N$�Ns'I�D��LԧM�PQ�!R5%&J�XB�?�@$�BaP�d6�D`�5�T��bQ��v= �E0̕ds�?$�d�]/�LfS9��m7�NgS���}?�PhT:%�G�RiT�e6�O�TjU:�V�W�VkU��v�_�XlU�m�����m�j�$�74�n�@����R-rƯ�I&��X<f7��drY<�W-��fsY��w=��htZ=&�M��YQ�{M�{m��w+��Q
�m���^3����2yN���ry\�g7���tz]>�W���v{]�.�X�[5-����<������i�!�������?_��������,�L��tЋ�׵ �,����nk�����J��������LUől]��eƑ�m��GB�\�4а96�R�"��A4� 4�?̥)ʒ��+�̵-˒�/�	�w�М���R#��îd>�8	�'��D�;���=ϓ��?�A�s#2��.���,9#��K�84�t�Д�5MӔ�=O�EQԔ�<M<�FC0ۑ6�s|C8�ӝ/;T��u]ו�}_��a؉�ODU2��r2�$"�]h)�ӭ�k�͵mۖ�o�Mc��T�VQ�}!7RV�+9D���yޗ��{���}ߕ��D�V]f��}#hҏ��:^W����%�☮-�����4`Ul�u�7n�u�1��NU��n]��X�)���d5���fY����Lf���.���L��.i5f�s�YI�-kiZε���
��L�%W�U�=`�j�����[������sjK���;n{jg�����O��ooz}т]Y�b_s�x���	'�=���/M��OUկ�]2	��e��sH���ړ���֪�s�'>Yt#�G�yO����o����a���E�wNՐm��|�x>����/���O��������ຟ�ws��m��������PN�����{��7���_�#4����(	���PnA���~/e�=�,�\��4�P���=�1�P�CR�,"i���9W�
`�����Ch��DI�Q.&p�_�;��E������[���&�ؽ�a�O2'å����7N �8# �Z��1�X���y�M2��$�L%�ОEw~hbċ��FH�#䄑XQ���8 �\���C�	����R�RJYL���	4.�h~�aTqxPV:Jym-