N�T{2N&�N�S-�Y+1\"$:y6q����\O!�[$pe#�v{&Ջ1�$�!
N���wPT�a%�b�s(w 7�#ag$�S#~�O1(W*/f'�n(�s	�3���"~v _`O��[Yf[/�[��'
N(_N�S>e*�!\OYe$�v�cY�eNN
�R/�S`2Ye2eg	�~2�%pe�g:NeQ
N�V}Y1 +N3N-AS&�[+�^Zf'�m*�s$�^\�_$  N*	N.�N5�Q20R'T8\8�b7o.�p8�v!�~7�8��8��1��9v�<��'��8
N �e*Zf%�l��*$�bR	N*N͋
\�S�Reg� :$
N/N6pN1ZP:T,'T,,T6�T/fU6�U8�V8Sb/~b5�dD8n@�s6w#Q;�:�:�
N2N�S;�S0,T8 _0>e+�e1/f&eg0�l>aw*��-����;ߏ2(�'<h��"FT�_$�s�w$�m0R�vb	�
N&ZP(&^.	g����.bN!�N`4/fw*$N�e"�l+��-m��yf[��$`N/\O.�S2�T;�V1f[?\A1\2b-�sB�v'T{+�~2e�>p�>v�Aэ>ߍ>��=��6�A��5K�.$$ $N0b0N0R�[/Lk/�v�/��$��$��5�+�7�&_4l$$	N�R
N8N,SO5\O:T/f[5�[3�_:`#b2Zf:;m1w9aw>�2�0��=�:��6��@	�:$DQ$$$$�T$$$$$$
N?�N@ZQIJU b9�eE$
N9$�S$"k $$�_5�$$AS0R&�S%�[�[&eg
T{(�#:Nx$${k�v��n ,T4�T/�['�[/r^/Sb7�d0>e4Ye.�s0�s;w*�7��7��7p�7��-ޘ4�*N"(Wb g#,{7�9r�� ,g1 M4 Rh K� I$ NB
NNL-N9KND�NT\O9�Q@�SM�SP,TJ�T<(WHYJ}YLf[6�[8\K1\HU\O8^W�^P _?U_Sb_V�`TaT@bOcc\�cK�cH,dFHeIYe�e6�eL�eO/fG!jMl<lY;m>KmRoL�oW�v,awO�w\�wQ�yF{<�~@�~J�Wh�R��Q��E��S��9��VۏKݏY̑0��[E�\�C�T:�T$���`N$"`NJfNSO/\O-tQ:�R<�SD�VB�W=f[#�[:\GYe.�e9�e7;m�s1u3�v2�w5�y&�~@�Fe�6��J����F�I��';�M�"$HN(}Y �v ��/��(�[[�)Y	�V3Y�e/}*��- wUf�uN+�PB�P(�Q>T1'T65TB�U9�V)Y&}Y%\7 _4�`4�e	g4�gB"k<�p<�p0�p9=r6�s3�u4<w>/}"�B��7��<��/��.�+�7(�4UO�[�Y	`NR)0R*XT/}Y0!h#u�v"�0�)�chQ�k�(WU_��$ N6
N,N:>N?ZP:wPC�QA�S:T=,T@ULfU=vVGPW=Y4}Y31\.�^C _:b?�e@	g;uL�v%w2wAGw?zzA�7��:��C��A��2̑&�7�4fb7��~$�v N<
N8N4N*O7�P3�QD�S2�S?�S=�S/�TC�V6�V7(W44Y>}Y/^H _1�_?�`+a@SbC�b<>e6�eK/ftfO	g4eg9QmK�p:�r>�sHw:aw3�{7�|H�~@�~B�O�A��;=�Fe�O��1��,ɉC��=��?p�?v�?��Kэ;ǏCُ*ߏA�7ޘH�Dl�J(�3:�<�s6q :y \ON�p�~D�g +s)��b�NV�vGW�eN�݋O"�Y\ �_%��0�� �eg�
T_�^ 6R&�S#�[(�n$�v�$N$Y}Y'\-�e/f1	g'}1/}-�~4�/��*��3�`^y!�0R'Y�p#��'�#{�&^��N�paw"�~��Ǐ%ߏ+HNO&/f	g �{+�~#9�<ߏ4(�/�PgR�Q�s�_-awɉ:N �R�~� N5
N=N,_N-�NO2tS=�S:�S<�S4(W(}Y7�[@1\E\:�]<�_:/f0�v(w5��B��(ߏF�F��(�5K�)
N �N:g��
N.�S'�S"�V+>e+�w��*N,Kb'c7�c*:g/Lr/t5u'�v,�w�x7�{,Ô,�#N$bT �4Y�$R)K{)�vX�y}Y$0RYe��	�v7�0RMR�~�0R�$0R��$
N-�v,{-�|2�%GPf[�g2�XT4f[�[$^
Pg"Hh2x9��!�O&f[h C$ N0
N>-N)?QC�Q00RC�S5T=TAT?�T<JU=1\<�]Cb?�cE�e9/f3 g