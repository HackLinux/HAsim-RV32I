Y�M��%���?Å�2�}���K�O��@�
EK�e�FӞb���YG/R����0n���;���'�Sf�ع�ޭK��&ߏ�`2�Ѣ��Қ$����A�>qH����ی�j���ℋ�s����hs���}�f�r�Έ�N'�!�ݧ�J�MYx��X��TG@>�x�D0�7��}��\�㒶W���Ť��FZ�j��&
$�e�Js�Zq���1e"e�|��HVd[��Z��H�k��BTf�����"��|�v�\��HՂ����Q���"�\�g��ɡ"���c��fd��Lm�Lq�I��V�Nüy�fjG3f����M���plj��ܬR��Ւ����5����6�]Y��JQ\�<�}��
�L��?c &�*Y&[O��f2�M}����kl��R�

��s2�',#��M�����E��]���G�"&�&x����Z�c��9*���WW��H)�޴�#�|�:��ˈ�6*��5�k�QJ�~Z-��m�(��Ns�ku�}-�?���� h��3�(��e�BDΰ����3�S��)�a��t�8����ǳ��	���kU��X	��� Ռ�0[���D�����X��!a���F���}�B��x#�}aa����-�"�X���*G�PE0_E��
��P͐������"��m���&{Gb��㻂�9#�i"�
� ڠߣ�g�ԍ��G8���.炸��"��v-�O��x:�wK��;��j��j���o�q�޸\��o����e�����(��@n>�{Q�NQ�XLٺ;�M��2�ҩ�A���o�4Y���M#S�m�q1�+2#�t��c|�$BR�!�ĢA�%�%�Ċ�b������:�˄���M�Z�h	�ã��0>�zT6\��o
o?�2�;{��y}�]YP����C�,�;$P&��q�-ܨ)}с�3���y�ҙ=Ф7[!sD��'�g���n>T��1�5�;�}Fy�&vi7>[
�t�}�w������@����J�tE`-��t��y%���d�K��9�eك�$��q�u�_$�����&�O��r^*�q��c����и����<�}#���ǁ�B��i��>גּ���f��g�w�^)���ɻ��b�ڥ���2��U^9��DR+��A�zEE�6��X�*�eB�*`�+��K_fugw5ʥ�q��� �T�Ѝ�Q���f��%��^���}�6(L��Qq;�I9©�2������e��j��ИB�q��h���1Y��
z&bX���%nX`�M���C��ᥝ;�$���&pYʱ�).� L�5G�b[�Jf���KeK�r k=r'��ɄU�)�s��7<�b#��D���w<�Ʀ�IwH�'���=�;�;��}'����}kI;`��6��=;�r��n�`ޞ�gG��B?�?��]~�E�e��N��΅�NlJ���t[5���-G�W�5*I?��q{��~�e�$�Z���$���� ���O$O��%ye;a;�s{�ڥ�
�͚1u��VA�� ���T��'�&����U����(	[�����e����C3ވ�A<F��<����VW��`��&���+��+�������.����r�6P� Q�.����B�2?f,<��e)�����ڄ��zg-)5��2���N̂�oq���j����T��	�Ae)�ج�� |Ff��[�����Ґ�I��r�1�SP女�%����%	�ŉ8�u�՚M�J0J�B���.$9ѹ��9�54����K�3ΛɟUT��C�a�ܖ*��x:e�F�$�#�I
,V��*QK֋�JҺ�y��F2xj�;�.n�s����=�Y��Ś	��`��3����MN�Q�Cيι�����C`"�	%�O%�}����ߤY�5b�ǌ+dHS`p*x'��?3L���P���X/�����B�e,�f�0��� �H�'��BBj[� $���Br_%�K�ӷ����fFe#�|��Eh�P
@�bϸҝ(f^wsҭ\?�F�1F��N�Y�W���.5k�>M1�:��z}�ۮ-q9���;2�)7�PL��iZ	K�\��LW����Q�<�(���� o~B!߭�X�������0)9q@�,�m����(��^��N)��/�t�sTP�Ez��#���T�RW����9��X.M�(�#�O�l��M�o�WZ���uyf��iQ�`����j��Ǡd��[�,���>�ݭ1��6�1��)`Pw�x��	�!#����{za�gwmQ`"���a��!�E�D����v�"L��r���G�W
QQ����hM��ç>N�}12d>8#�c14��c�C�f�Y&C���C�&��
ͫ ݨ���"t#��tH�Q�؝��w&Ǽ�¯�T���Jm�F���(+CMM��21'�_x����>�,/�XR!���1��a�M��ȟ.7.;[,4����~[��-z�* ��9Oj�0�7~�z����P�»d
@v�pj��"(��<����P�yoӈ 	)��Ln|	^t�g@�bC6��Ժ�C�:�ZƸ�op.�ϵ����᰹���L�{`��̊g�k1����k�8�(�pD����w�(��	צ܁�Gے����֢yU�E:\Lr�Aڮp�A�@�g��p���%fJ��EH�ƍ�2�Y�1��Rb��f)�^�X|���]hb�-F���Q@�#��=��4F��>��9����&ك����F��=�,������c�vÚ�ӭ��|���̴>����d{V�C�4f��.���jUһ��ޤ�0_SI�H���%e�0;�p3�)�������=-�{"����٧���4�������٢���fo����I���ɑ}�3�����A�U	���6W��lt_��hI(�� �H��?��l�,��L$E��_ 
-ȓ�=�`o�e��"S���VO���3$'��/����<�� �Q��Wy�)���:���	�|�D�u�4��ߦ�$Ч�����@z��1js��G%����'C=c�l��b��y	{cb��������"�$����
�p���т ��#I��H�����_y����mI������Y���4�e-9$���m���@�p �U��H6J��gUZ���R�j�֮iWɻ��=���&���%#��iN�3Sｏ9�<?s�cp�C�)ɵ�\�%l�'�;
}����p����V����OT���Rq�8��AR��I-�h�����+B��Q�)S��tRA.��8���ڌ��0<��L��"ٽ��aߤ֤`)$z	Z-�m3.k�C��2ٍ>N��s��H��ji�Xp�Ҏ�OLֹh=�L{�l�J�"[-���%�bg�~Ë��x��@٭gUj5���;��f���̗/���V�➃�0�[�C"���d32�'��I���ŕj��8˯���%��x��dd��1\�3{�oh����'�v_k�3.���q{(��~��M*n��FH#�$:<�/G1�t �׎��Z1H�Y��f
_�x���A��I�	������o�̟���D�|�Tx�u6"�Mi�l�d�
���C��d�9�Ok1Mӡ����[���C���5
R�Q��"TQ�P�t[�|�&�g�(�������ڄ�yT�r�x\V��[�~�>:���E��E9l��2	oG*��j�\F˙(L۪(k�:[@t1�V�E�2�"��U14H��S�Lp]@�H�:�ĪLoy`�5$�6$!T0�H��L;p����Z��/���5��z$��җ{�i��m>㊲�"�-�g����MN��y���a�:Ӳb.~X����~O�dD��_�<�jO�:�;��)펰HW�E��E�-�t~��	�8�q����/�_���2�kY%M�H5��v�
i\4=(��S�]r�ưo�=�������k���d� r�������~�b�66�-�Z�ׯ��T-�EQ���+v��x}$M�f�����WC�	'"RȆ��dEc/��Fdc���������;�ق�~+>e93�މRȇɫ���?�n�U_��h~�����̪�G���ͅ'�.�A�����2�挕8����[��e��a���SUT2)��sl���Ϲ:e70�b�"�Yu��sW�,��td�~O��D�x*��"�T��G�NT�G�=d+���u�x�K���|SU�H!�˺jȨΈ���B�h)��I{�h-H�"�����Ck��/%=S�ͣ��a9�i�._���/re��W��q~���p�{�|S�q�g�}�;�I���{���$ ��n���?�@�Os)3�d�