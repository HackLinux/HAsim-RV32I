I[��t��x��C�d��	{����P�PϪ�"���3ܥ����B���[��M}vmm��
��z_;�P=y�zӫxea��	��޿�
f�`�6���,����TO�%g�/Y鳋�,E���+1P�#��¬}v�s���*q!Y)-IJ���G�k�c�L[s/���8����죑�}�z':�@O{/mb��i�zg�	mL�y�0K}�Mw]N�Ŀ����*� �ӨS����4��d���ME�y%�]�-�r�Z/~���}G��s��>d[�Cȱ<�d(�3����F�2Y��T�}7xa�`\b�N%hrFD��$��H]9�ǉYLp%\�I"�h��yB�����H��'{�G���اb~���bz����PY��u�6��L����,Xz����Kg�&���e|�*ҥ�)BT�O��w��Q����;�A'�/��C 4+���N��;I~���sM͆�b�VM�6�)��l �B�X��%�sY��ॶo�b��c ��6>�2��tk<��.	m��]/^J�=���+�������e���D�]}�/�n�*���i����{y�'�<�_���q(�2���4ɾ�x��A�n��������+���yKD}��Ի����+��]lN�m��[���P���Y��RS�L��h�!R�����*y1�a��C�<P�S5�&%]l�LU�k�!;����u��hj�v�Mb����ju�5+��*.};����g�1���h�?�I�;�O<��.G  �C�,�����'�y�j^:�� ԫkhxp0&G����)1G"����E�/y����xU�:|亦>.�is�\�6�>	��ߟ#$sݴI�m9��i��O��W�B7��m�ꑭ��(G��R��9v� �~2��9z�&@O��JH�����0�Op�
�4 �B7��G.P�V���?P�S������B�F���J$��>&�k�0��f4jQ��?���|u����2�c�| e��r���쭾)�?���b����������?�P�K�2i}a��<�4������#��&Z.�`�fJ9����uK�z���l�O<�ŵ?�co����|�3��A,F��/5���-�V����xSm������,����\� ɯ�/���y��J�gy��¯^�^���?�W:�ָ���8�G���p����)m���|7w7���l��*�y�.:�c1J.�$~g,�څ�W�y���{�.��<1}T�q�8���z�E�ՎZ��ߘ�/���ϊ;G���m��9�%��?�yt9�MnO�YH���e��E������Mmu/ ���Xγ��[� �ӯ��,�Cti�׫��?���W�&` ������^�i�H��*��m�������\��'�E�z#N)�O7�����9�)����|v�y�� S�Eb�|���f~�e�p��~>�t�	����P37(u�;	oKl�=
މyJ�P7G��V̇��K�����f��^��B���һ�8+RV���{���e��TܼV�����W�P�/��'��\l�U����J�`�쩆	� ��8G�l����;,��j,(�����(�`�n�^��6�T!S�Rؕ�{��mx���f��s��m�f/�ʚ��p\d����u�_�YS�X��e5�G4�Y���N�
A��m
�c����sBb���P���	����*�O�5�x�:o��GC�yR�*�F��p�Be
-��	H� ;���[�F��;|�;�Q/�)˅���jTO�!�<"?1�&�:#��*]���)x�74��N��x�!�����U�DJ����+���Z(���v>�l��G�2�y����M��Q�(W��|
�i!���y0&�g�
L�r�L��0ڡ�wܣ�O�{� ��z���	�����s��Ϟno��Z�X������^�Z�����zf��]aw,��G��@�Z^���B���B���V��Q-na����g�Oý=y�2?�'�E�0����AD�%����SP�Q����=,�f����t���#j�)�GO8���N�"�w���K��7I��7���Z����Q�?���.]p�ފ�H1{���|݀��{i0`o�q�9<������Cֈ����N��Q�d�����=(F��7fP/\�PGu�]���%Y7G�U��j�x�<mo����5����+l��CӶ[�E��M;�w񼙚��ؤ1s�M���ФϦS��5jٰD�,T���ڪ���mґ��I_�M�Ԧ�,(�41�Ф���YԜk�9�ap���m��8m���S�$���4jc��Jz,��l������Ctm4�ژ�k�7m�S�ƹfC������"dV�0�.<�M���k{1[��z���>�n��~�O98���^�V�;2�h��w�����Mb����������l�sp�T����e_ڛ^��w{��s}r3�H�7=�?Θ��Oq�S0��-�L���N���ke߹2��{�FFpJ�|](mp	�����0%
�ص�d4�]�2�щ�"\��a_F/��3v�hI��2�?���ڠ&���#�p�^����Fmx�zd�'�"�x[}��=5�S�������g]"��-A�\����x�EK燝�lt_擦2��yO�E�`��{y���(,�$1mR|�i@F��YQ��ȃ,�`��!0,�1����[u�!4p�~&���pH�d�1��w���q��%n��_׻��5)�Zm
�,��(��8��]�*��T�9"l�$�YР��p~H�������?"W3O������_�����gо�V0�1q��mƯ7�i�C�h�xD�<����ֿ��u����'�����0�]y�\�,��țP���=qIw4K
�>�lv�D�w�"�f?|�u98��>Ǟ�w<)��\�M�zA�v%+���vSB�W�^�Acݩ��^���j�+k�#�5���G��~m������k\��	��P��]�30����%8�n���;K���I���z���/�r��p�mq���n �/jGZ&Ο�:�L�����6���uHC�]?���(����'�,V�'�)v�tj�Oݣ��_^�#<c�x�����/����������9�I�蠁�U)�7ӴG�l9翠R�l�4��d��C?A}v&�zD���0��7�`O��*��������,J��q,��/'{,� �[]ެ-�J�G����%�x|��$���LD�}��i�f�M�DI�ʒ��������(f�͎J�8����ڮ<:�2�W%�+�f(�Θ�#aI���Hy'`6`IB,�QT4BPA��0�娣�ݧ�s��xns�f_K�Aܰb�e���{��mU�0������w������;8M킏�H�.�`�a~�'�N�^/����F�G���"}i�Q �E���4ӽ��� ?]�\�3��F2�	���;�[Ǔ?���HH�<%�-$�m$/��f���=;�;Try���r$0��	o�	��O�p)%�q�K#�	�������6uh��Ť��7<���?�=�5����~q�MQ��.#���i��!��b�"�?�.�OcoĈx�F</��.	�lb�v�8�в�PS�Ԋ�0?ޟ��Ԧ�C�}���C��j�N��p>a��t�U]_t��ћ