                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           < K  ��� ��� ��� ���    �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ���� ��� ��� ��� ��� ���    �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���� ��� ���    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ���    �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������22������@@������������������   ����    �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������		��  ��������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������YY��  ��77����������������@@��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������..��������������������YY��II��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������11��  ��������������������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������cc��  ��MM����������������������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������

��--������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������nn����JJ��������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������jj����SS����������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������AA��  ��##������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������,,����������  ����''��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@@��..��..��..��..��..��22��HH��������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��������������  ��  ������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ������  ��  ��  ��  ��������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ������  ��  ��  ��  ��������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ��  ��  ��  ��  ��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ��  ��  ������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ����������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������