������Ѳ���uw]`��yk����{|nuzzaez�|ho��ohtssnnikv��oi���ov~�}|xt��}{xy~�fZVm������ɹ�����{qx��p����z�qynogknmvglrxqhjlldhomnrzvqtysomnqfULL�ڮ����ڨ����vjZ���az���wziw��nYs�~dbrvrgiidmungiupqilonqtynlql`O�ư����ڲ������h���ys��{jiw��fq��gfsof`dbdeorpilrnddnjjdkgQR�֦����Ѵ������l��������{{rmuu{jzxkbldjdb__jgrgdgolZa`jjb]Nj�ɞ����մ�����}s������}���imx~{mrowrqiU^fnYPenkdi`YdbbWVWPY�Σ����γ������w����������wdw��qjmmmge\Ycg^\[\bgd]_XY^TJJ\��������λ������|���������upun|�p`lpfhfWR^c^UV^jj^YXXVa\Gf�������ˮ�����������������vty��oeeogjd]\UfdYYYY[`UQ[ZSVMc��������û����������������oqr�|nfaacslXNS\\eaSPT^aYIHTZ��������ι�����������������rw�qig]cmqf\YU[ZZ_\UV\ZOMX[_��������ƶ��������������}��}{�{klrh`eic^ZZ^]VWd`TU_]V\ZM[���������������������������~rv�vmvtabja[_YS[XU_dUPZXQ[_Qc��������Ǫ�������������~sz��}ytfmvmjiZP_fXW_ZW]]Y\]UTZQSw���������ŵ�������wz�����st����rdhonqraUZ]afbXV\[]fbWRWW]��������ǹ���������~����xqt|���|qpuuqoica``ccbbdgggdegdec^gy������������������������~zxz|||wqqw{wxvlioojppkjljinqnmmknrlrzz~��������������������������|w{|wx~zv{�wxslpuvsswmlmprxvonopuytvtt�����������������������������}~~{y�uzzrotrsvunsoqxqswmqspptxtvy{~y|�������������������������������z}{{yzzyyvytpuotrswsrsssvrqsuwxzu{x{�}�����������������������������~|y{||w{{xwprtuywqrwvwvttvyzxvoy{z|�~{{�������������������������������~}}{z}|z{{ywwywyyxtysv�yywm|w{|qu|u~}y~y~|}��������������������������������~�~x{|{{zvzxzvxuqtvyrzxwxrxv|�s}yxy��}���������������������������}���~�{}�{|~xw{}y|zuwzpx}utxpllwt}�utmz��~�ty�~����������������������������}}�x||}��{{wsr�zsyosrovwutqlvzutxps�zu{wq���������������������������������~��}~�yz|~txpnsrrylipsuwtzmnymz}xtsp{|~zyv~����������������������������~�~��}�yuwyxqpommplsojljxypnwtronpowtpuusz�������������������������������{y}zz|wolqpfknkkmpnhmnmqtnpninps{qiortz~}���������������������������~|~����zwvrmmihihcejifggdknijnmijllprstqim��������������������������~xz��~{yytmkjea`aceffhiighilnnjjnonkinonlio�����������������������������~z��}vompnhhhdbcdgjhddfefkmnppoqtmddiouvonz����������������������������~��{xwsnpmfda^ahigffehkjiiijmrrqqpnonkmpqrttru�����������������������������{xyyyyuojiigee`^^bfikhefjmpurlksxzvnknssrqty{z|������������������������z|��~y~�|yw{|uhekngc]^beccgfbejoonmquvtx|ztppswxtzytz���������������������������uz|��}wxxz�xplkilhd^bdhijfeinmjkmptwxz{ywwzyurty}y~��}���}uu���zz������������������yu{{|�toy��|rghrrjgb_`gjgdcckpqpqsw~�{xz~}xvy{}���~~����z�|z~�xsx����������������������zuz�~tszzzyvopohgllfdddgjfempkkrtu~�~x}����wt}�}}�{}~���yu���{ts{�}svzvv�����������������������v{���}~}wtzvlijkmmd]djihhfdjqsvwsqw��~|tx��zuvw|��vy����zx��~v�}~�~zz||z�����������������������wxwwwwusrrrnijpphhjhfghjhiklosvwy~|~��~|{{|}����{~���{w~���~��������zz|z����������������������~y�qsqpwulkoqkrrffmqlggbfnopompx~{yz~��~}���z����yz~~��z���������z~����z{��}��xz������������������������~}�tkqyqlmokqrnigosojkjimsqmnvvwwy{{~��{|����}~�����������������������|�����������~����tx����z�����������������|~~xrvouvtrnqt{utxrs~qtynqzwnx{sy}yx|zy�{~s��t~�xx���t��u�����z�}��v���}�y�|�|�����z�~��t��v��t��y�}z��s��q��{}y��{q�yu�yu�{x�s|�z~�zz��t�x|�u�h��g��i~�px�o|�n�~r�w��o�w��s���t�r|�u��u��y��p�|����k�o��h��k��o��a��f�wy�{��|�w�~z��~�v����|�z��r�v�o�}s�p��o�h��}�zx�v|�h�}r��~|�w���~w�x{�l�|t�q��x�~��q�x�p�x{�y{�u�x��u�y��j�}�o�zq�ry�v��y��x���l�p��u�~}���|����y�w�}�q�y�t�i�}�y�wz�n�e��r�r~�}�~x�{�u��j��n��k�tu��s��V�ux�l�v�t�{|�z�k�s�z�v�m�q��k�{�t�q��z�t�m�u|t�j��n}�s��zv�g�~t�c�g�xt�u��w�p�s��s��p�sz�h�s��t�s�t��o�p�}u�q�~�~z�|�s�f��v��}�r��p�~z��z�y��r�zx��s�}s�m��w��s�l�v��s�n�}y�^�r{��v�p�f��y���y~�|v�l�v���v�q�{y�p�p�r��{�t�b�f��o�\�\��b�U�s��t��x�z{�t�v��p�]�oz�o�s�x�~}�y��u�{�k�i�{y~�d�g�|~�y�y�w�����s��p�uz�q�m�h�l�v����{�{�z�t�x{�p�x|��q�h�p�p�p�s��b�l{�n�l�`�y~�u�p�n�m��l�|u�i��r�o��x�w�q�w�t�r�r��i�t|�k�yu�d�z{�X�\��q�z��t�n~�j�q�y�z�s�s�u�o�x��}�s�`�sx�g�su�P�`��X�e��e�T�]�{u�v�z��m�r�}��{�s�q���n�p�q�w�x��y�}��z�x�v��l�m�e�o���z�n�i�z}�f�q��}|�~v�r��}�|�v�w�q�|��w�u�{�z�i�u��y�o�h�~u�g�a��n�b�{t�c�x}��p�v{�l�l��r�s��v�b�{q�n�|{�v�t�}{�p�ww�f�xu�q�~x�r�m�s����w�s��o�g�~�q�w�u�q�g�c�m�u�w�z�u�~y�x�w�p�y�s�v�t�u�y�~�{��y�o�y}�}{�~��y�||�h�n�x�j�z|�~x�z��y�u�v|�{~��u�y{�q�s�x�}�y�|}�z�x�~��v�s�u�v�w�}�v�}�t����w��z�x��u�~z��m�r��y~�|�y}�k�xy�w���x�w��u��t�{z�t��x��}}�r�|�~�x��s�s�x~�z�}�x��q�z�u��v�{|�x�v�i�x|�~�~�o�rz�t�e�q�r�k��