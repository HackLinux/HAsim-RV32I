w��医�l5E����9��ͱ�I�UQSu�t=���c+<=C�{��TZ���օ�L6��9S�����3�)q�~q��t�k�&����ΌPPvw����*j�;Ί���VE!/�B�d|���1�Ԁ�y�ƴ'=Ksʓ�%/*�ͫό�>3L���ڸ���k�y���+\$�J,��kqk>S,m<��d���Mk�5A�5����E7�Z+Z٢V�z�wԢ�鉎��髿D]�xј��1�b%W��%O�[Wк�S�_������}e-�З�b��y+�Wv_�KJ��o��y�bu�k�W%u�u�D��$��(��D��|5�0}���Mŵ��A�.��t�œ�ŻH��K�����AKϖM{ҵd�M�,Z���V��ܕ�Wګ�����Wk�TړE�{=�9Vu	�E��i8�춢�h�&�,���x���j�hn�Fu-�5���
���������޽��Vy_�9Oԧ�~�/�އ�ܧ=�*�]*�]N:����ͼ�V�#�ݜ*M�jQ��¥��;RR=[q>�����ꆫ���}��'����o�lS�>N��f]��欪bgEW��J��]}*E���Z:�!|O!2�����ތ�qo��yo��p5����?^͔>_uv��
��.�%Q���.�j����L�s��=�Δ<���s�j2tvd��=2��1G��ͮ���y�����F毞dd6�$#�񓌌�8�,dmasʓ�!m���n���E(��g�?�3�Bs$���u]�	_;%�Ϻ����>�v��	��5�b/H�{A"�O>_�~�p���
y�%����G�Zh�T(��{2�)���Z<Y0�
�6�cYg�ZP����u咎\R�b��vd��cz�1}O1����.�M{ ���OљB�9��/=���O2���,�*�^i=͵�-�#�7�K��N�b'
J���(^*ῖ�X��{��"=���۹ų%#nZ���V��Z� ����UБE�{��*���>�o6�USh���}��?�Ny�]���K��������Q�����D�u�[A�����p3�)�p��6X�}�Ż\�jv�n���d.W|4�����r��aλ;�9��9��0��4�B��iaEt����#���X�|^�%=-�;�\��U�.<�/<�o)�|-���ŷ򵔬|-��:[J��l)��-�5�ſ&����-�/[J�ul�}�������������8����h)�����ˊ_,_��%�����ſeh)�3��6-%����mC��������_�ZJ������_�ZJW�߲�R�n��,\-�\-H~Ks[�w��?��Ҽ�䢤26���,���c�F*����)�_*ɇ2ag��4�꼵�w�YȻ/&x/�����fzT�R_}���^X�Н�U
6�|x�k�+�#�7��J�_��b'|��%|WJ/��_�Y�\Ž�^���W��]����iO+X��;�������qs^d�^9�hq�PX�н�*_xY"�{["_x]"�{_"��P����&�ܠ�/ _,˻��w��K��[y������@�{q _xs ��/�r>��������~?��A������+�������{�|}:��ͱf<c����_���_~�o��A��N��]d�{H�;�|�aj��45��j�{�|�:��,�8�7��|
��o�(�#J��6_��ͧ�Nj��%�﷕pnD����&��˗���ջ��y�r������6���N?_��罽~����v���v?����K6�yo���m���n=�ۮ�[�oo�/lW��j>��4��o�gK,�^�ɻ��!cΧ�tqq�{C����mz�]M���Y\	!!Bu�����q7 �CK�]	X��Nj�� uA{�Z��*���âh]T�je� �!��j]AA�U�j�}E�DQQqE)U�[�Z+��d��ai��������m�g��M�I2�L���@qf����x^���ý�4�����:���J��f��<��"7�������CwO_��B��[�� �u��V1�^��=/��3��y��y��P쉐3`�Rz�bA�d�!���yɖx�ѐ���3q�ӛ�\�<��`E��++$��ȾR�Q>�Q�fd���Q>z�}�4q$��0_�����2T�<C�!	���A��rk)g�����`�����|�g�A�@�@э@��@���u��{�zTz�y�+����������!��C\_���qM�j:�ut�+�^;��j�������ݗu$e��M�}�'�����{1`�n";��XYC�� r�f����kyh��G��)7x��3f,k
3����<�*1l�!�I�y!�膊^�+�C�9�ɭ����tO�}הīU���T������=��0���>�SVD*=��7Z5f��U��7��9�g"�6�����e�����1�6�V�y4R��4(L_���Lǡ pږX�ʁ���M )v�?)�pP��I����J:}:�]������Y��N/�:P;�WN)����J8�@p��������\ ���Fby쥞��Ѡ_�����0���~�7�|Ï�n){mi�w��|;��[DTa��f���r˷>��>��gSGwl��Q�a�L �}�;�{Q �X����$o ��t��t��������=�e�}(Z�ܴ�"��l ������|ŏ`Y�`��ؒ�)o��߈7Y�S:���ǹȏ+�p���
��Z9�6�^�� ��x@��<��\�1�
� �v�&���7n�9p�<�+
o|?��W��9p5��<����#�.����L���go�p5�2�F���U�~�{�W�������������2p۩	|��2 ��VMzգW-��ߣW]���B\]��Y��Қ��@�F��mc�o�݁k�[��{ ��	�e�B�|���O����P��H ]��0�'B���(x�g#��	��A��@z�����o3�j�G�����dT��Q�Z����\��=<�&z�L�����B׋�3��g°�����0�n��φ6�~����Q��ƌu��(��}���%ҢZ����!/�6�	���$|�����q	
���%�*c�Oߐ����+�QP ���k�R������ѭ���W�H���ui��j4!R~���_�RX��.!ʝZD7i�n��t�����"^ȕ�}i��Cy[*�Q�Wb�c|i�b<�yżPY�ulSXyG���~nFy�
|U������*|y^�GT�+��U���0Ov����5� tz����Ų2����5���if��e�r:~G[1��P��o�]��+h�A��\�7��;��[�{2 9����ש���{z�Q���Q�䀯��<�Qط�>P0����!����������2y=B/VnG�qŊ��?��`�UU����r������W�2δ/�<ބ(�e�#e��w�Ogo�����/E��/��.\
800 ���P ������	`#@#����k "�W�,,,���r�G�� �L���h( ֩Qy<��_ų��8;��K/g8��f�N�,�z���4csz���|_8[R�bh7�.��1kS*ۙ^C��K���M[]]GQ	�pv����������>l��@n�1��Z݄��)G�)��'L�ucḟrΘf\&�Kb�|��]�:!w�붷�/��$LY�e]����1���X��D��"9 ����x�lЇ��cEKxpe�6��ɣ��^�,�h�U��e��׽|�y�u��7sw�&~l�ި���mF7����y���g~<+ꬭg�����b���0��gӺ����'솎�*