������������PVFCR70(4DKlz����������������VIIC>3((33Rdz����������������IF627+(&(7Rdz����������������II-1.#&3Cdz����������������IQ-1.#+Rdzz����������������FB61.#3J^zz����������������FV-5>)#(7Wdvz����������������IVI;C.+(3>Wdv�����������������VVI'JWC.37>^pz�����������������j_]8-^WC73KRlv�������������������zojjdW@77Rlvz��������������������zzzdfRRWlv����������������������vddpvz����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ucc�����������coy�������������u�u��������������ooo������������B!1ET����������e$5NH|���������eFE:Hr���������eFbAHm���������q]ROAr���������kFTOHm���������eInaMb���������wITOSr���������w_~SSn���������o]bOH~���������}_ZSOm���������qPrSMm���������kInHMg���������ePZHMS���������e]RD=`v��������eQC?3N|��������eV>3+Dp��������_<.(&2j��������o617v��������eF5+#Rvz�������qV'Z>7Rz���������zz^@Rv������������v�z��������������������������������������������������o������u������;^�����F7|���|_%:�����],A�|���e,/|����j,/|����i,/||���i,4x����P%3Z����I#E����],.Z�����v^����������������j���$���6n��Bb��6Y��;1���|� ��������{��{��s�{s�{k{{ks{c{sk{sc�ccsscssZ{kcksc{kZksZskcskZ�ZZskR�ZRkkZscZscR�RRkcZkcR�RRccZsZZccR�gg{RR�JJcZRsRJ�BBZZR�BB�BJsJJ�BBkJJZRJ{BB~: �99sBBsB9�99�91kBBZJB{99RJJ�11{91cBBRJB�1)s99�11s91�1)ZB9k99{11k91RBB�)){1)RB9c99s11JBB�))s1)�)!JB9Z99k11{))k1){)!R99c11R91s))c1)�!!s)!J99Z11J91k)){!!k)!B99R11B91c))s!!c)!J19J11991Z))k!!k!B11R))B1)c!!R)!c!911J))91)Z!!111B))11)R!!9)1c9))J!!9)!J!B!)1))B!!1)!B!9!))))9!!�  9!1!!B!{  B)!!9!s  9!!!1!k  !!1)!c  9)9Z  1!1R  )J  B  9                                                                                                                                                                                                                                                                         generic46    2          (   (  (  h    