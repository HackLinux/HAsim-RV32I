�U��B�EċMċ�U��E��E싍����Q�U��E��E���M��U�E�+E����@�����A�х�tP�E�;E|�F�MQ�M�������E��U��B�E��M�U��D
���}�E�M�ȉM��U��R�M��T��뎋E�M؈�U�E܉B�M�Q�M���R���E��M�� �E��UЃ��U��E�   �E� �M��j���E�M�d�    ��]� ���U����M��E��H�M��U��U�EP�M��y� P�MQ�U��M��P�E��M��Q�U�E�E�M�Q�M��K� P�U��M��P��|� h�  h��* h8�* h�* �:� ��蜐 �E���]� ���U��j�h#�' d�    Pd�%    ��  �������E�   �E����������   ��i���E�
�������   �E��E��E�
�M��o���E�	���������   �i���E����������   �Th���E����������   �/]���E���������t�]���E���������d�����E���������D�)\���E���������4��Y���E���������(�� ����E��E��� ����X���E����������O$ �E� �������B������������������������ tj���������������������
ǅ����    �E��������������������E�   �E������������������������������������ tj��������������P�������
ǅ����    �M�d�    ��]����������U��j�h�1' d�    Pd�%    ��$�M��E�    �E������MЃ�������M�d�    ��]������������U���d�M��E�E��M�Q�U�E�E��M+M����A�����B��tV�M+M���A�����B��t<�M���U��E+E����@�����A�х�tj�E�P�MQ�UR�EP�M��"O����]� ������������U��j�h��' d�    Pd�%    Q���   SVW�e���4����E�����}� v�E܉�0����
ǅ0���   ��0���;Ms��4��������  ��4����z uǅ,���    ���4�����4����P+Q����,�����,���;E��  �M��Q�� ���E��E�    �U�RQ�ĉe�E���4����Q�U��E��M��Q�ԉe��U���4����H�M��U��E����4����T�����M�Q腂 ��j j �� �E�������4����z uǅ(���    ���4�����4����P+Q����(�����(����E苍4����y ��   ��4����B��D�����4����Q��@�����D�����L�����@�����H�����V�����W�����H�����P������P�������P�����P���;�L���t�ዅ4�����4����P+Q����<�����4����H��8�����8���R聁 ���E�M����4����P�M�U�ʋ�4����A��4����E�B�M�d�    _^[��]� ���������������U���D�MċEăx u	�E�    ��MċUċA+B���E��Măy u	�E�    ��UċEċJ+H���M��U�;U�sD�EċH�M�U�U��E��E��M�Q�U�R�EPj�M�Q�������   ���E�MĉA�%�URQ�e�EċH�M�U�E��M�Q�M��  ��]� ��������U����M��E��M��U�    �E��M�;tC�U���E�M�M��}� t(�M�� H���   ����t�E�P�� ���M��M���E�    �U��E���E���]� ��������U����M��E��@    �M��A    �U��B    �E��@    �E���]���������U���$�M܋M��  ��]������������U����M�E�H�M�3҃}� ����uR�M�Q�U��E�H���U�J�E�M�P;Qw
�E��@    �M�Q���E�P�M�y u
�U��B    ��]���������U���   V��l�����l����@��l���A3ҹ   ���u$��l����B����l���9Awj��l����  ��l����B��l���A�E��U��U���l����H;M�w��l����E�+B�E���l����Q�E��<� u �   ��Q聈 ����l����J�U�����l����H�E�3Ҿ   �����E����p�����p�����t�����t��� t-�U��t����
��J�H�J�H�R�P��t�����h����
ǅh���    ��l����Q����l����P^��]� �������U���,�M܋E܃x u	�E�    ��M܋U܋A+B���E؃}� u	�E�    ��M܋Q�U�E�E��M+M����MԋUԉU��EPjQ�e�M�U��M���  �E܋H�M�U�U��E��M����U��E�M���E��]� �������������U���   ��d����E�����}� v�E���`����
ǅ`���   ��d�����`���+Q;Us��d�����  ��d����H��M��}�s�E�   �U;U�s<�E�����}� v�E܉�\����
ǅ\���   ��\���+M���d���9Jw�E��E��d����Q�U���d����HM�M؋U���R�V� ���E��E��M����U�E�EЋ�d����Q��d����H���Ű�d����H�U����EȊMֈM׊U�R��d���P�M�Q�U�R�E�P��������E�M�;M��   �U�U���d����H�U����E���d����Q�U��EƈEǊM�Q��d���R�E�P�M�Q�U�R�������E��E�    �E�E��M��M��U�R��d���P�M�Q�U+U�R�E�P� ���E�    �M��M��U��U��E�P��d���Q�U�R�E�P�M�Q�� ����   �U�U���d����H�U���E���d����Q�U��E��E��M�Q��d���R�E�P�M�Q�U�R��������E��E���d����Q�E����M���d����B�M���U��E��E��M�Q��d���R�E�P�M�Q�U�R�������E��E�    �E�E��M��M��U�R��d���P�M�Q�UR�E�P� ����d����Q��d����H����t�����d����H�U�����p�����~����������p�����x������x�������x�����x���;�t���t�ዕd����B��l�����d����Q��h�����h���P�y ����d����U��Q��d����HM��d����J��]� ��U���$�M܋E܋H�M�3҃}� ����u
�M��
  �݋M܋Q�U��}� v&�E����E��M܋Q�E����M�U�R�y ���ԋE܋H�M�U܋B�E��M�Q��x ���U��B    �E��@    ��]����������U����M�E��M��U�+E��E��M�Q�B;E�w�M�Q�E�+B�E��M�Q�B�M����U������]�������������U��j�h��' d�    Pd�%    Q��D  SVW�e��������E��P�M�U싅�����x uǅ����    ��������������A+B���������������M�} u�  �E�����}� v�U��������
ǅ����   �������x uǅ����    ��������������A+B��������������+�����;Ms�����������  �������z uǅ����    ��������������P+Q��������������E9E���  ǅ@��������@��� v��@����������
ǅ����   �U��ꋅ����+�;E�sǅ����    ��M���U�щ������������E䋍�����y uǅ����    ��������������J+H��������������U9U�s?�������x uǅ����    ��������������A+B��������������M�M�U���R�s� ���E܋E܉E��E�    �M�QQ�ԉeԉ�<�����<����M�Q�ԉeЉ�4����������H��8�����4�����8���������������������������M��U��������"�����#�����#���Q������R�E�P�MQ�����R�������E�M����U��E�PQ�̉ẻ�����������B����������������Q�ĉeȉ����������U������������`�E��������M܉��������������������������������������������������;�����t��E�P��t ��j j ��� �E������������y uǅ����    ��������������J+H���������U������U�������x ��   �������Q�������������H���������������������������������������������������������������������������;�����t�ዕ�����������J+H���������������B������������Q��s ���U�E܍Ћ������J�E�M܍��������P�������U܉Q�Q  �������H�������������UċE�+E��;E�  �M�U��PQ�̉e��������������B�������������������Q�ĉe��������������U�������������E�   �������H�������������U��E�+E���M+ȉ������������B������������������������������������P������Q�U�R������P������Q�������r�������B�M�ȉ������������������M�U�ʉ��������������������������������������������������;�����t��j j �?� �E������������B�M�ȋ������P�������Q�������������E���p�����|����U���E�+�������|������������t�����x�����x����U����t�������t�����t���+�p������A�����B��t�M�U싅t�����P��  �������Q��l�����l����E؋������QRQ�ĉe���h�����h����U؉Q�ĉe���`����M���U�+щ�d�����`�����d����������������������������������B��������4�����4����E؉��������,����U���E�+�0�����,�����0������������(�����(����U��������'���������������������������� �����������������������������������������������+� ������A�����B��t6�� ������� ������������������� �����P��������P몋������M��������������E�M����������������������������������������M����������������������+��������@�����A�х�t�E�M싕������J뾋M�d�    _^[��]� ��������U����M��E��H�M�3҃}� ����uR�M��Q�E��H�T
��U��E��E��M��Q;U�w�E��M�+H�M��U��B���M��A�U��z u
�E��@    ��]���������U��j�h��' d�    Pd�%    ��   ��`���j �M��� h~+ ��q ��Ph~+ �M��ל���E�    �E�P�M��4x���E��E�X/( �E� hT�- �M�Q�O� �M�d�    ��]����������U��j�h#�' d�    Pd�%    ��l�M�h`�3 �E�P�<v ������r ��t�,jch�, h��* �M�Q�v �����Az P�v| ���� jT��w ���E��E�    �}� t%�U�R�M��b����E��E�� h�* �E� �M�M���E�    �U��U��E������E��M�d�    ��]�����U���X�M�h`�3 �E�P�u �����5r ��t�,jch�, h��* �M�Q�\u �����y P�{ ���.� �U�R�M��!   hd�- �E�P��� ��]����������������U��j�hH�' d�    Pd�%    ��t�M��EP�M��v����E�    �M��h�* �E������E��M�d�    ��]� ������������U��j�h#�' d�    Pd�%    ��l�M�h,�3 �E�P�t �����@q ��t�,jzh�, h\�* �M�Q�gt �����x P��z ���9� jT�=v ���E��E�    �}� t%�U�R�M�貓���E��E�� t�* �E� �M�M���E�    �U��U��E������E��M�d�    ��]�����U���X�M�h,�3 �E�P��s �����p ��t�,jzh�, h\�* �M�Q�s ������w P�z ���~� �U�R�M��!   h �- �E�P�K� ��]����������������U��j�hH�' d�    Pd�%    ��t�M��EP�M��ƒ���E�    �M��t�* �E������E��M�d�    ��]� ������������U��j�h#�' d�    Pd�%    ��l�M�h��3 �E�P��r �����o ��t�/h�  h�, h(�* �M�Q�r ������v P�y ��膀 jT�t ���E��E�    �}� t%�U�R�M�������E��E�� �z* �E� �M�M���E�    �U��U��E������E��M�d�    ��]��U���X�M�h��3 �E�P�!r ������n ��t�/h�  h�, h(�* �M�Q��q �����#v P�Xx ���� �U�R�M��   h܋- �E�P蘸 ��]�������������U��j�hH�' d�    Pd�%    ��t�M��EP�M������E�    �M���z* �E������E��M�d�    ��]� ������������U��j�h`�' d�    Pd�%    ��`�M�j �M��x� hf) �>l ��Phf) �M��=����E�    j j j�E�P�M��$� �E�j�M��6� �M���z* �E������E��M�d�    ��]������U��j�h#�' d�    Pd�%    ��l�M�hԌ3 �E�P�p �����Pm ��t�,j@h�* hܛ* �M�Q�wp �����t P��v ���I~ jT�Mr ���E��E�    �}� t%�U�R�M�����E��E�� �z* �E� �M�M���E�    �U��U��E������E��M�d�    ��]�����U���X�M�hԌ3 �E�P��o �����l ��t�,j@h�* hܛ* �M�Q�o ������s P�v ���} �U�R�M��!   h��- �E�P�[� ��]����������������U��j�hH�' d�    Pd�%    ��t�M��EP�M��֎���E�    �M���z* �E������E��M�d�    ��]� ������������U��j�hW�' d�    Pd�%    ���   ��4�����4���P��( �E�    j h���j ��4����������E�j h���j ��4�����$�����E���4����A0    ��4����B4    ��4����@8 ��4����A<    �E�������4����M�d�    ��]�������U��j�h��' d�    Pd�%    ���M��E�   �E�E��E��M�M�U�R��( �E��E�x0 u�M�y4 u�U��B8��u�M�y< u� h�   h��* hH�* h8�* �Ct ���{ �E��M��i����E��M��$������E� �M��������E������U�R��( �M�d�    ��]�������������U��j�hh�' d�    Pd�%    ���M܋E܉E��E��M�M�U�R��( �E�    �E��H8��u	�U܃z< v$�E܋H4���U܉J4�M������M܃�������E܋H0���U܉J0�E������M�苉���M�d�    ��]��������������U��j�hh�' d�    Pd�%    ���M��E��E��E��M�M�U�R��( �E�    �E��x0 v� h�   h��* h �* h�* ��r ���Gz �M��Q8��u� h�   h��* h��* h�* �r ���z �E��H0���U��J0�E��x0 u,�M��y< v#�U��B8�E��H<���U��J<j�M���$�%����E������M�膈���M�d�    ��]���������U��j�hh�' d�    Pd�%    ���M܋E܉E��E��M�M�U�R��( �E�    �E܃x0 u�M��Q8��u	�E��@8�"�M܋Q<���E܉P<�M�������M܃�$�����E������M������M�d�    ��]������U��j�hh�' d�    Pd�%    ���M܋E܉E��E��M�M�U�R��( �E�    �E��H8��t� h  h��* hؚ* hȚ* �2q ���x �U܃z0 u� h  h��* h��* h��* �q ���zx �E��@8 �M܃y4 v*�U܋B4P�M܃������M܋U܋B4�A0�M��A4    �,�U܃z< v#�E��@8�M܋Q<���E܉P<j�M܃�$�c����E������M��Ć���M�d�    ��]�������U��Q�M��E�� �~* ��]�������������U��Q�M��E�� �~* �M����t�U�R�a ���E���]� �U��j�h�' d�    Pd�%    ���  ��?3 3E�E쉍(���������P襓 ���E��}� uij ��l���謮 ������Q�pd ��P������R��l����j����E�    ������P������Qj ��l���R�������A� h��- ������P�د ��(����M�d�    �M�3M�_� ��]��U��j�h��' d�    Pd�%    Q��  ��?3 3E�E�SVW�e��������E�    ������P��~ ���E�}� t�hK  h��* h��* ��n ���s ��ڕ ��E������M�d�    �M�3M�ĩ _^[��]����U��Q�M��E���o�����]������������U��Q�M��E���������]������������U��Q�M��EP�MQ��f ����]� ���U��Q�M��EP�[ ����]� �������U��Q�M��EP�MQ�:� ����]� ���U��Q�M��EP�UW ����]� �������U��Q�M��EP�[T ����]� �������U��Q�M��EP�MQ�UR�EP�ZD ����]� �����������U��Q�M��EP��A ����]� �������U��Q�M��EP�MQ�UR�EP�" ����]� �����������U��Q�M��EP� ����]� �������U��Q�M��EP�MQ�L� ����]� ���U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�D
 �� ��]�  �����������U��Q�M��EP�MQ�UR�EP�MQ�UR� ����]� ���U��Q�M��EP�_� ����]� �������U��Q�M��EP�MQ�UR�EP��� ����]� �����������U��Q�M��EP�MQ�UR�n� ����]� ���������������U��Q�M��EP�MQ�UR��� ����]� ���������������U��Q�M��EP�MQ�UR�U� ����]� ���������������U��Q�M��EP�MQ�}� ����]� ���U��Q�M��EP�MQ�UR�� ����]� ���������������U��Q�M��EP�MQ�UR�EP��� ����]� �����������U��Q�M��EP�MQ�UR��� ����]� ���������������U��Q�M��EP�MQ�UR�o� ����]� ���������������U��Q�M��EP�MQ�UR�� ����]� ���������������U��Q�M��EP�MQ�UR�EP�s� ����]� �����������U��Q�M��EP�� ����]� �������U��Q�M��EP�MQ�UR�E