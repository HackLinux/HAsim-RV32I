��x����
   ��x���f�@�3��x���f�A����x���f�B]担x���f�@
斋�x���f�A(���x���f�BM���x���f�@|؋�x���f�A�E��x���f�Bo܋�x���f�@����t���ǁ�   ��P ��t���ǂ�   ��P ��t���ǀ�   0�P ��   �v�   �o�M�Q�&  ���U�R�EP�MQ�&  ���U�R�E�P��'  ���M�Qj��t�����R��t������   �у��E��}� t�   ���t����KTCE3��M�3�� �����]ÍI �xP EvP �vP �wP ������������U���$�E�E��} t�MQ��:  ���E��}� t�E��  �} u
�  �  �U�R�EP�d  ����t
�   �q  �M;M�s
�   �_  �} u
�  �O  �} tN�} u�} v�  �3  �6�} t0�U�R�EP�0  ����t
�   �  �M;M�s
�  ��  �} t�U�R�EP��1  ����t
�   ��  �M�Q�U�}� t�}�t���
�  �  �E�x t
�  �  �} t/�M��U�}� |�}�~��E�ǀ     �
�  �j  �} t0�M�Q�U��}� |�}�~��E�ǀ     �
�	  �4  �} u�M�ǁ      �U�ǂ      ��E��M��  �U��E��  �M�Q�U܃}� t�}�t �<�E��P�M�QRj�E�P��/  ���(�M��Q�U�BPj�M�Q�/  ���
�   �   �} t(�U����0  R�EP�M�Q�U�BP�Ѓ���t�   �o�} t8�M�Q�U����  