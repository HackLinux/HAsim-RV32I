�8â�PU�������m�sK���]w������)���:h��Sh#���]�̢=�F�X�_�G���3���\�%X����T�!�:��^�X�/T�����3�|/�3�s�ZZ�r{�GE ��d
���sQ�3.���0���xu�C��z�ȭ�#�}:�����,�u��=��c�ʖQTө�����z�p�PQ�KxR����窸�=.a�@I�˵h��r��κY'�<��f��t�jcۻ�yn�=�R��RT��i��������_~�3H�%��c�hc-�/�0i�������ȅ,\���
_�(�a�g��߇�?H�S��^Ї��+�-��~�	w��~Yc��_Grg����t������¤-��t�u��4��X��Np\%��4*��ٶ�".��y��<��
i�(F��וD)%��!溠�7g��`�O{4s�r�0E|JQX��`ʬÓEr��:%��׉������ܤ��Mt�AP�At��!�*D�[RB{UhD�T!��=˖�ki�j�N*��=ԧ��TjU\i��S�-��>.�C=pLH�'w��븢�k��m��)�|Ü\�?ޜk.��d�5����\Ϳ,���;E�_��
�9)�҇���<j3��-�;�� ��;�d����%rx����6�r�����(~�^[��HSj|}�Y������a�w?�h��%H��׏Dk�p��ߤ�>�v2h$5���b�=]o�+�90zC�0�f}��M�a�&���A�qO��;$��~����,�ƹ��}N�����Ob$=�z#�-n���+����n�f�T�� �����t�*����C�.F/��Ɣ_z���a���C_��g�B�
�Ƥ�������>���1V�k���Y	Y�D�+·�NdE���59�;
�ű��=&�]֯����*
�Yf��1d�(�P*��e|�q�33�W���g��ηA��-��3@F/:��Qۉ�<�;Fwnu�������@TyX �D�7U�7H:��3��^�&ٱ�_�̯��Z�U�O�^�?l����C�ۙ�@W���E�_���2����I��.�'MҔ�v�(qigf�I���~�L��k�?i<\dLXY����`��5����,c��^�NƷz<�V2|A���?���1->R��j)$��^ѢI'����JYO��E��VROh�{,&
&��`�=��V��L��&����՟+���a���:}��1�9"����0�L��i�����S���zrϘ���1���;:9���n�tb6ۯǤ�h&� _{7�\�w��W����@��"�&���x���k�����g��+Ή�[�0�{�ay�01x���_���o ���k~�������/k����d��~Y�N���hf��'z��?R�	k�����.g;�>���S�=�J_"��c���X3!�Z5XB�{\�y<�Χ?K��6��u�ɢ�e��w����q[o@�_aȢ����'j��1����5ƦU@N�X���(VH%���͖Tv�L��1m�W��a�2,u)��S�6�*[/���}��i�-/�� �G��QEҒD0��|%x87��i���r���L�����e��� -�JR�"�:ק�,���K1�|,�q���>�Ɋ�i��5N��6�pj�N��jC�������������ŵJZ�L8.!O�EP�TE��6�cw)P�]W��x*]B�(�Y���r�c#ze�ޓE���gj�A����`퀓�*� �j����.����M4���u��8�B�,>��
��ۃ��f�%�A�F�v�=�*���9����}|�^��-Ɨ�#+@�?���|L��0�|U���v�e�=}�@�T�lg��{�����bݖ卆!_��k̯&�z��<�؊d��"��>?�T�W��8�Q�K{�݊V���\����֑aЫ��_���7U]���}��	�B���0h�E
�ZL��mӧ��ڴI��V�X��
$�J�Ŵ��%�~C���Ca�(*�':-}�e������+*:� �|�ܗ/�����;y��{���;��w�=gt��~3��K����_��5��KΔ�Kv�ͷ�F�U�Ş�$_�*��_��{��|��I
�6SaD�X!U�_>\E��k�����B�g�&$�D�@�*_9�`j�3;�P��%Q6J��kt�{F���7�T{����ڐ�[��B��
m�B�(	^@�-�F�����?_��O����>�7��������_�ݹ_��K�y8{A�������{�Ǥ�V(���r��r�X��:,O�wD�޵QN�Krwݗ1��=��r�ۃY�r��R=�1�;$w����'���|%��qN�n;S�1����1��!����{�h�r�����9���rw�z9�'���w]�i�y���]^?�쓂�,�kWx��7��5*ۧF��]qK�i�^�fx�^�{≋��,�q�&��B֩q���/�+��}�4�oD�	�vOG�<�`���jg�H�	ٙ�f$^�=����?B뗪�����&wK%�4Ģ!��S��Gam;��a�lA�%�W])PJ;g����- ��'U���Mqa%*�aU��"�4�S˙zc@.@���,���.}�F�[���W\L��J$؁xX:M���5�d�ToԨ���7Hh�������h ����3��	�j�ő?���t�T���+<���*���ޤ������E����x�?�9��2������t��&MKJDd(��Ձ@ �$,���թ_"w��{b���tO�y&��qnƑn�H��ޡ7e��r&���st�T�S��U����O%sͱ���X�cf$�҃]�}���ݶ"ט�E���Tڬ9N��=������O{_P��Ւ΁�gw��w����b��X ��/xQ�����C�ngB�n�FПZ������q�No�Q�x��
�C:<3��ܹ��3�]Wq������ATdD&�N�Å�H W���Ԇ¯�s�2�V��kP��D�Ԧ���}�FW�(�UE�a4[E�(�*�o�o�}7�Meb����$�]�&[��'"7P�HQ
���I��JTQ͙xE�C#yh6n�%�G�%�)�p��~����a{s���'��~�m�����1�{����#S�?�>j��;�G����#͠�l>�<<�u_�Ѹ{~r�>8�Dr�0��+'x��~L���+5�����m�P��E�2�W�}��6�^��ܲ��-�_پ{�>,6�b#g}�iw����+$���c�x`�];�M<Kg=�xv��mٴ���9��w�Ev�Uɷ'jI*�mWN�i2��+SO����5��>w��7���<+���7�JS��>��^e<�@���0|��fR�@�g��w&��.Ƴ�up:�Y"��Kds:pQ�x-��ȹ��ĩ��7]��q��^����=�}FG��P3�����=Pa�gN���3�q�}�?��q�W4����\m9U�𧲨3)�U�rm5���8��`�q�i{�H��9�~�z����. w�Ƹ��#f�����5qJ�V1&���|M�ʕJnӘXt�����Tٲ�{*�xװ�Dن߿KʰCyK�|-�~UR�-a�Mgjʼ�ݎ��˰�8�XRY�-��{�A��u��hͼ�y���nZ���Ty@<4�^�3h�A��v��)�Xz�Π�t���XCg_�B��{<�*p�j�f�w�m4|ܯ2]p����K�����~��K Ƹ� ��S��F1��*�@� ׿�)8 �#�� �" �_D���ũ��/���b�N�>������ ���H�Tx-h%S0@+�6@��g�J��V���J� �J.�: !b-�X�vty:|؎���	%zI��8#4G��p,�g���1�ޠ��E#����$5s��< #����A���x�v`�ӕg�D��\TS�i�[RU���Uy*U�3øY��c��ص&N��'�:�s�@�z��F���4���JÍ�4��J$��Rb��eq���4|w�}?=��GKR" �%5�,�<�jmh\��>�7�-
�'~�p{^8����w�����j��=���,&�Rʓ0e���t�!�dcڿ��|���ޠ�;lG.��-f�{�P1� g��{��J�%�	�=�FOќ�͖Ɔp*��娟�/G���Ї.[������ M�/�$���']eA��u;�	�I�a�>R
��:�1�7vT� �6���;@�=Ҹ��^�d?��@Dɖ�ɡ]���mȩ7�Yu�!χ�נ�p�*9C	�i]�_��9��f�ҩ������N:�=aj�O;E���?�&
���w�w����x��n �Dߏ����`��3$
����)Q����Mb>��Zg;��lt��c]��&�uw�%Q�3����D�������:����x;�zl�(0e�G��o�0����B��Z���i9��82��1�r�7 ҟ>��(|��Q(�O3�hYA<�m�w�(��>#
8��G�_s��r�z$}�,�����x!F�3/
�Cg����K^;yaM������g��Gj��'��El����D���8 >!M;�Z �_^����W^�Rw��"�7��Qk�p��m���ɿF���@�ч7W����7��E�|[ct&A��mNl۶m[�|c;L<�&�m۶��o��{NW�����WW�fe�Ѻ.ψ�����	�25��"F�_D)+�F�R������ ��uE� 2�%
x���.C?���|{�.��z��^�������c+Lp+��N73����[�N��� ���m*�>������WRn�۹�
L~�;A���R8�a��R��b�'J$�^��O�xѾ���
h��~�p=�[-��KO��_�8׾&����0ע�=HW��a��}��V~��Z*@�˭>�tg�#WIL}���J��uЧ�>ٳ���[Z"#4�LeDt�n�Ӳӷj���.�Ar��P��V�<�Wf���-����s�r�)m�BP����:����򙷗H���#�u�g�Q������Z�N��ۤ*�����-g���`�c�����qlѴ��-L}<�iB(�يt�h�3o�SZeqz�WXawQ�����d\QJ󗐧�^P����e{��Y_3Q��(b�4�H��Hv`?��6I!�;�"���|��z�ӂ���1��G�`a�mk��S������	�A���qi��4r:�e�[�T�;>�D�q8$P��R4�2v���m�
������M�/S��4�Ǚͭh��q�k)�����z6v��o����!�����"�5���x(��_j�4�-!�l��r*V|��*�m�لѭ�W*����`P�l�z��DXa�i��7���߻����������&�0�H���$�v���������r���!¯zj����^\ë{p@n�����C���~�u�77�d��'�SV�}�����J!�0.�w������o���0�� ���T�.E���[�)�YY�<��/C��`F�]�e��`p]v�W�#xA��ܕ���pf���O�̇�1%b��텚��-���Z���v�j�*����pJ�;haU�޳�t�<��MO#6��Bs���k_�z��1��g{H�"0���:�N�Ӈ����:�|�����zHZ����y��v�I�>*�ј��j��HV@����u,�q�ѯ�g�Q�Wid԰�^�p��S��	���3�R��~څ�B;�v��!�y˱~7�W��i�yi���sFv�l������$E_Z���m�-�l��u@t��C`���.H���;{ءѓ3�펃P�v��}��͈J�X��+Y���r�b�'+Q��g�?�����/�'�'�����x�
�6a�=^�sҫ3?�Y��)KMl2r���(�
д���2�N����鼃�z)��ݹ�����[y��&�cp8��˕����mV��pè`;��g��AP�,��m>'pi������1�݁�.�ӥ�,�e�Ì��l�m���B�9��"99/ѫ�ɨwp\\ȴI��e*�ؚ�w<�;�c5���~TC@�aƞ������(��U���H}��Uc~F�)����s!���� �� ��u���Q�� �AX<_Pn9 �"�)g�j&��G����={0��T��m����L�>o�|ـ�_��;�ut�څ�{[�E��ښW��1�U�����:w1�I��)-b7��ن��ڗ�%B����C�P���$�J���i��Iu]}�|�l�A)a�:=$e��鉧^x�E��}i!�ӟ��QPC/���/3 ���	:Qa��+�z�߫�DV2z
R���b�3���z'S&��t�l�s6Ф7&�
<�\��(f��J�	;ܘ�����7�+�� }�} n�8H(>��.u�s�K���D�H�d�3[/ ����1����z����W'�1)�0��EK�OX�� d����l�,y��F�@�������E�l6Ҭ����يu�,�ܐO��� ��	�5� D ِ�D�&��d�d�b��f��r�=OJ��+r���fp~�[��d~�Y����SBz�G���w�o�)(Y
�z�LR}���"ڧ�7���	z���g*��堡b�ml;����S�;�� ��!����=��О�RE��b��j�/5|�n�����T}y�6�6cp���̕چ����{|+xO���F������Z���F#�L�v$��vn���g���Aݞ*:�Hy�a�APj0<`�\�g\r��4��I�5������
֘�U>��P������>8���;�x>��u��s����?h�ϻ�iFG�\b�'T}�q�ޒɕ�TV{^47�GT����3F���'Qc�[������W��&�o�VI��|�vW{~UZ�~�l R0a�!�� ���J��In�p�MnNﶒ�6j$��x/8��Z��[��J�\�ƺ"~��_Ɏ�R��L�����oF6AH+��g� �����<μ��!�Y~�SC�Ȱ$(���BF�L>�U�K佊��Z}��t�T�X81^�����*��2�$�F�jY>w��X����V�f�hM�tꠍ_�<3�)�$Z�f���.��w1��ˠ�+GQ�4��C#cs
��� �S�0;�W�=�p���4�r#������t\�4�OsĐ�j�����5�+��<&"N����TY��-��n�,ɭ��~{���N�Q�f�nQr��K[z������}�x
����OK���2%�M٫���+h��f�������+d��)3"���1k$�%Ѥ+~Jm;+:n,���U��O���@wĺ�;�j뢢i�rW�[�E_�s�ک�]r�k ���ܤ �i��>���/1ʞ��uc/������d���J��=:�Ѕ{w��x'��j���v��э8�v�=Vo_ʠi����۹b��ݬ�Nޝ	�T�ѫ#[�Qӎ�t�S�Y�]�(�Zq��Vy�:Zr�R�=�E�;�a���
�n��`$��7�+���{褊��8Gƛ�\j4��d�d� �G̒RJ	�|�<s����I�|��<�E�����Ϡ2�uw^�C�i��Y-��	����dU�E�5o�kJ]l�Ŭ͉��+���8���m2�0O:^:��ܶ;��ݨpq�k4h:�\���
�3�J�T&�J��NcONu.~(]9q���7��MfDk���őmR��u�P�+9U���`��H0i������C��k�=o� 9����r,�N�A�j1��êUM�ʯ��sLM�v~�e즒4G���.ٹȔ��໪CpD^�Q�yQ`�����u��'���D#��_�8�\��oZ$K�|��Ý��g!��6o=%G���s�'���6īZh�T4&�}ɀ/���J\����6o�'��Mk�����K�mN����D�o��J��P��ʨRa�^EX29w5���s�<g��e��A�J�B��a�Rw�����3Ǭ�d�����f��g�����Uc��M�
�=���WO�ɜyS�.��06�;�
�Q@|�[�^�玑C=к�"F�7�+�k�������F�J���I�&�8$�Yz����=� �I��'�.~��~�q��0�0�R�&=\�h��ȟ�e�(�?X���c�&���Ra�f�֯������Of[\�HA�J��,'h��hT���J�_�<QU.�\����!�Y\��
�O�J��y/��V�x�oc�k��ʣ���B����RxH�Mlԏ�@68��΁,|p�2�� MI�c{
�V8���;~-p���5FJr~���ˑ����N�%�_8�v0Hħ^��/	�3�2�2�҄�! ����
W	�*߳��%����X�����4��'#�]�Ծ��<2)��Tf	�΂/��E"205������7x��3�]Q]*��<�D/gb��H�q�;/ư^XgDc��-��	�gvX͸F��Si���4R,ۻdE3�x�����6�n�͔5ί�����n�i��a-��rx��'+j'� ��o��o���8�c�7����^���C=G4�L,�|�F��o�db-��$�p�|�q�F��?�3�)oYάJ�/y%���9'��L�:?���f�����HJ�g���\��M�n�Ӏh�#����g�����R��ž�9���/��<��$����I[��&���1�T��@��FѺU��F팩J�����]b��-A�*�� 1������*���
g4&�����_L����-��iCtF�;i̯ƽ�b�C�ڡg�C��/�����a�t+u�]��7	$��~�n9�7eKT�	���
���Ƹ�A��J;��YO���Y�����ݻN+��	���k!�����9_"l��)2qAy�P�I��1�0����<���������?�4��T�ez�����\���d�Ԭ�3�
�|��o�����/%��a�a�����S��� p�Kz/:z�.�S(���3��ҏ3z��9�ɚW<ɔ �N�oe���&4�`�4�s���#�[7�?b��I�U��9E�G�t����y����/���_4�-�㿫c��>�"qX���0u�
`�D�|���Z3��O)�[�l�F3#�6b��VA[��|*,׮;��Z��y�	����M:��15�sX�����6���N�v�v좆��T����5;�K�ZwW�!�)��,PF�M��&q�L$�e�������]�Y�59�������Y���h����i����[���Jr��ms�pY������.�y�b�:׹ ���k�vNr"`l$ϒ�cJ���!
��Y�4H�8�M�>_-�;G����.�A`��l�E���]��]�Ǐ���HfL�E����ٲ�4���Å=���@�M1)L9��L\����,Z�)�}�s�[�.��������퉆��S{|.o������wO~R�;u���~VE_�7r쉢��d��?��*K�F'���$����Um+B~%�c�r�K���I�8�T��hK�7������l�%P�.�ϕ�:C�Tz�r_I�ʭ[.�^��BZ���]��Hj�����쎔g�Kq�-pR~`p��������{!�s�'��|�����y^+Ʌ`\ڢx��Z��s�&x��a�.2G�ݜ�,�'$��x�����io������t�Qh��p<��]LB�#w�]��'8nD���^���c
�Ǆ��yMq��;��ȟ�ad}����7	h>q��w�����,l/�]=k�x�>t�Er��t�U����.�zH
#rW��]ٽ��KmWݤ?"�)3�}�	UP�.�����Li3��=��G��S���ˁ2ɲ�FxЈ����%����sk�vV1�o�D��wV��(9s�u~���x��6`�s
|'���@@����>���b�}�n'�h����i�v�Z�t�@%C�g�9's�Ԁヿ��Qȸr�����O���=�����e�v����06��:?�������XaN�_@�u��������4��ˠ� 5`�p��筈� '<���U0�"4���֌ד}KS�d�|E�	����$N��a{��ɣ��PS���i�o5O(���k�h�<�`���.9���E�!��T8k�I� ���GwK�|�����u$��������/����k������)��"C�Vdt6�]o�pϩ׬�s��DL��,"����qaZ�Tsw�Yz����"~����d������P,��		�H�=�;]t�`�����+���ŷ&�fa�i�~-Ů����-i>�\̢����&$��-�HD��9�4�2o�"3�ߟџkJȈנ�:M�i]�'�y. Oa+]_���C��]8lx����p�g��KD�.��%����H4���F��=���'xo,=	�Yׯ��	���%�����S��u������|�B��ZѾ�Vt���=ҷG�=��YvӾd���c