�����N �.Mq�/٥������q��>�PrT�����
��Q����𲥏���K��C.�*��h��Ss!�1n���H�Ղ���������E33��;twU���ѣB�&��>����.{��º�A�����-�5��f�V�e]�����M��xY$%F'��.s;�u��=���8���c�(ɋ�i�K�N+gH�mga�����Z|
<i�����y�/o�2P�@vذ;�t�ބ�=v}X��lX���\�[0W�mhZ�M=��P�oU�S���xtt� J=��-�FOA"�%J�'5�>�-ڟ#�vg&넉Y�	�-����#��w����p��I���O�!T��mfx����%vF+'tc����n��G�~�Q�԰�ֹ�n�b�rp���~���Y���c��+����}IC��o�����N�|��9��K���o���(��^oR""u�Y#�N��s��_!Wsoͧ'�T:Ct�\�\���u�%�����K��kJbx�>��#�ޒ�ė��ks��gdM��U?ﱿ�F���DX�Qˈ���nVf�4r�)�&.�[�i�K2�+��,()���jF V�-G��w��q�6���lm�2�C��LOU1^"���BAK@����Ve���r@��Q�{�98[?nB����˯�����jY��W��]_,D�*�$*��@��m�=]�$,�	�x��ȧT*&�8-ے:Y��:����O�Ϛ`�,}���=��!ţ�<��)����qN @ �f@]ap-)sß�mN�_,y�i�=��i�B�9��X�\���H���?Xqr��*u��A�Ӌs��{Rq����
���I<��O�:��J�U�`sd�m�9�~/U��ȓe8�,����s������L������$=Alo0�l~/��q�7D�K��3�N�;���|Y��i�e�et0 ���)G�����ܼߣ��BXP���Z�ԼKh�	�qJ�����.|���^���%��B�bJ�Q�2K��|�g��I{���	�)fUV�}��� �6o�m�����J���[2V"�\s���2A6v�G�E�I�e�V�����*<h#@�=�*b�����Ɍ��B?X��v�0�_"ϡ�~�S�%�\h���5J��vhS5�Ŕ{�������-�t�O�n+Y�N/b�d)�[�b�?��!��G�
��Kp�0��H>S"+W�+�x�T��V�u�m!�|��GAM5U�7��~�½ ���hw+�� Po[ɵ��R�7��AA�}U<��+��n
�9A����۱���^����7�f)����ٳ���۩r��pۍ����W���aVր�a!�L̓q��'��>�r�|��v
2�;�˗�f�%����ᔯ�Q+�ˈ���Ć�m�+t_m�]~���Aqd����4�b���j�/;���w��Tn��J/5]n���������:�*p�����#[2e���v�C�HS�U�'�%�ˌ�^m���P��E�p� �r�6C�Oeo��_j������z��&��&�$8�8���w���9i
��dJ����pW����5�S�:�*��zi�)������?f�d+�8E��L�W��Mqt�0Q�p`������w���7Q�&�D�إ�g�� ��]�I]�~ձ!�׆Ɗ����B��g���5"YM��ߛѸ8��l���E	8�G���j`_x�zA�!��f��`����+�0���1K��ڰ{��@,$�Ƥ�1R�uX�0����Z�Tc sK?)���� �W%ޡ���*rV���,��e��y��)/�B�W�|�0`��E'U�V�[�"ؤ����o;�DR?�d��aK�pt0 aAIo
���N�����=&�;��\ �Y����;��HI˱
�vS\�$���P��Dpz�i����+)t	׭���)��YG���O㽟��;�z �A�X�x��S���3q�Ә;ўi�%+Rm'1�3���f����0�tXˬp9�z>@�?�)�(� ��3
`LӲ\!�������ɇO\�7�|���TMq���L�)�G*���nR�S�f;d�ah��3UNH�P2�(;>��3�I>zv�E��6lQ1�h>�	1�ĺ�Ŀ�[%�~����:�5�n ������'mQ_>����T��aɰE�,"s"�����"]�_ӳ�WΔK���bĀ'�f�D��3ªd���8I��m]�R�S�44��;�6ې���.I�V����}9@P�����k�o�[en���A\�fS�ϡ��j�Á�H�k]�0R�*
`D�N/��얇vJ};�Y#C�\I]3���`'�������WN"���#� e���:�����AW����q�PJ������[�����0Tw��g-r�T�|�����(3�z4��-����⊉��q׽j�-Gv�+c+��́������K�$M�Ս�d𽸦՞23�)9*�X�J�	r�(
�":My�Ϻf��nu�n�%Yd�3-��C����BpJ3a����0Ј�e�ݽ�;�R-��)i0b���h�X�D�>��5&�౾uW��N����}�1>z��1�-J�'�f�K&�Nį��m��.�M��4Z`U뱀�Q�VI3�I}�Sz�P~����a����
���&:�Ճ��-�<PF��6�)i�w&�?J >�T�o0�]-Y�?��H�I�{ߺ����Dq�Ŵ��K%1�@\R 4��n�p�O�s���]��:<a3�u�t��۹���ʼ�	~�i�-�x�f��w\VY����;��>&�)�ׇ Ze����#@��􄵙D�S��L{#��7��	����u���h��j�O��mq`uZ�V@��9xs�D�6��z�+Ç����Y*֋=��l�Ƌ`7wĢ��������L�ȣ�����,C(���J$�+��5]9�W�)RvW��mb�M��I��8c|g�������m���X;��GQ�S����A}�>g��Ẽ�kL@��m���\q�����CHr^����(��1��A[W�+0�~��x!>�e
�2WfK�Mp�L���݊N܄���ث��$������(�\҇�T���>_a�OĒ4]fl��7t�U�)���.����\cs۝4=��'9 Zd	��h�x<��:�1��a�\�$���|���961���P���/B,e=rM$���A9ڇ�u��QP�!�X�K��O��m�-�ϣ=�?��H�V�h�V���nmis��I2(s�?�
�5�>���M��Ru͹��k��(����#q�3x;�?���G�L]�+��ڐ�U�Է�y�R��M�$��6o�*+�p����쭐5uR��jJ�:�?	���M�-�y�j��N���Wc��oݑG�;��y��+{X��z�mj�g�x��=�/r�P���ʬ�F���F��vSц��!����W\���?�o��gv�.�i���%�0RR��A>����2�op+�i�>��.�(Ĕ����;{�9����n�S-�]@�
�R�h����8�vgz� ��f & wk�^-u��6`.;�K�1b��Ļ<����t�֭w�=����ɖmT6��BgJ}�}��}�{�� =�X�a�n-Z�B�0PI������/��~��@�SD�|T�[�E�U�5":�2����#�y����i��T!�9��牐����!}?�/��A2u6*������Q����f�(O�7�y���鿼H� W|��e4#���F�
�zMXZ�OJ��G�<�/�7�ǰ��*éC��(`K��!x����n�d$��M�w��ؕ�b�Ps��W��l�d��u���o��� ٥�(��e��6��K+�2��M�2�i�x����vG4�Wż�
B������.�H�Ȓ�1�K���"�e��<����!"|�g30?��:K���Y�H����#��h�Q]�����Jr;��WZu�?P%�K\}r�O��Ȼ��Q��j�u�1 D3��ƶ�2,�2�MyS_c[�N\4�p�i���p�إA���H:��g�>uY�Sţ�f�BN�Es�3��meR߭��6�)�/���ryK���(C ���«�ᾟF�$����ט��e2��H��s����^9ΥK��"�u����32��o�+���ꮼx�`���7�+iO�79�~̞HI����W?Y�E �����aC��sw�YC 3��t�QԚ���n�H%"����ѕ~	Z|����n{_;U���B.7,�),J�&��}:�~d�B>�t�bq����q�hISzr������e�r?D��LX����6�@zy=�-�Xa�Ag���ʷ�f�sd�L.�;��0"�񡹢�V�7���PKM`�^�i � PK   :\|A               META-INF/ECLIPSE_.SF��I��^�>8�k���rP�\��UZAA�V�у =~�BO��C��ֿ&y<f�[���D�J�Vݔ޿u���,��A���)������-Zi�/��_�q��z�2~�0ަXx�C:������/����s�M�������œ⿨�̳Ҫ����?xx��&꺌�������A�E�d���qg ��"�Ԇ���������ee xN�4��W�V�^Uu���Y)�����W����I�������Nkaj���M!�����Tr�2�״�:�Eu�U O���G?���;pqDvBv?-�=42}B�P��D��<�0++�m�������(�[�z,�������	'@�.��t	�w��c~]��ze^	��m��4o��g�5��A�do��)=O=S0|��EB�y��J�����m/uB#�[��x��<�H���3�I�C�U�sI�B/hҮ֡��嬲�d����������gC1\+�1K�F�0�lu�X���>$-��|;���H8�MK���Ww-E:���
����������W�"�]�HibTx��eԅ1s5W�c�[~�J��gM�Z%�k0gA1��!W�
����=߂J=��k|ʀ�4A��� ��ӏ��m�* �L����E�翟��Y�ï٠0tt�n�7�Mg]��5+FOEQ=�zs��y�*kaP0^ꕣ�J�����]{��v�]p�VΜ��C��=�9n?���pޕTz�W�=nɯ��a�yi�T��e{�Tf��}���Q�Z��pV�]ڍ�Κn_%'�^��6��鰕��[�b
*5n���C�u�5@��&�j�C��*���j]�,KH��5~h���<���@��t��q�l$�s��(������乙SPλv,9QK��v���K:_�Q�F��Y�x��l�q3.�c��r�_�a���х3c���~l��ͯ��DQ�4~a3^l�s�pX�鹹B*�°�9�?.�%�F%�} �E�!tGA�e�2G�?�Så�����?�W͠�ٻ}�ܢ]��J�^�
�^/Z7��>�Ay�����}VG~�</��k��3\�����sP*7��aS�C2�=�Ď����M}ӵ��"D��cE����]H�tMny����c����|3��y� ���b����c��U��ٍ�	=<�LΉ<�;[w-�f�;û���=b�����(5h=�^��dm�:R�ֻ���dW�p�C3��M�(�J}7	�KE�á^�w�?��uI�����hәВ�4P��07��,��_%�J��SD��/�λ�C��I�,��� �_Z�����'�����(/�__�e���z����̂�����O������^�i
��Ǟ:e�R�2�l2@\��	�0j��I#����W9e��6��0���VPW;h�'����H�\����S+@}�ʻ \+u�Y	��m@��x�	����^�?�Nժ��V��A��E�V�h���fa$�}I��	M��9��A�J�+'��.���a�y���B꠹wfs��p��� �K�7��&��vtP'y��;ú�h�s�K�ܭ�}z����x�P`3���q|���U���sM���MJ��w��,�@�X��2u��1���`8ltw/HJ��
��@^q��z�-�X��V��S?r�|����c
��Y7=1`����4����zI�����7��7x�S��[��b��hΝ�������$N��ۑ��W�*_���,Q�?�ѳy	툞�K?�`_u�i�>��qE�^A���
=sB��.d]B�9K=������PBOp*}����Px�b��~�ݲ{�ƍ֜�H�>G>c_ҧ�VZ�?��g�ް�KG3�VХS�h��-$�z=�Q�A����7 NZ��
�����(o�K�A˽eQ�������F $y �ԵJ��<et�*ó6�!�;՝�*�Kg$���֦�L@�������o��-�EC8?u�� �զ03=�X�2��M�Ė�<�������=�@�;�_
5'�y����}��k�zɀ���,�G:bC�����m���p#��"p���)����@��X������c���t��"�����~�.��x��XNo�V����X��
k�u�z͡~�.��"σۄ�c�Y[y�7#@���4y����x	X7��Z;��ap5T���u� T�~\7�����/�������f'��k��ú��9W{侩�M�V0�/�zv�b�t^�%ɭ�8\@o�����m�������;*Qz//|�iq�Z�� <��@��n�/x\A�kV+~S���ӈ.W�n/���zm��\/+��(�(�ߣ������F�Ы�ᚽo��:[gPP"�)}�e��]��f7�t���+�������$ܪ��h�+���W�>zβE7�`̼��*�����SL�se���K�v������ҧ������X��Bωn��i{�^ȿM�^���d/�w�)���� �sT�þHV���n&#���r5��P]e��..s��;���?^?3������%ɔ˵G	���U^Rl����l#3涃��%�>����>�Rn��̦�ޭYa�MeDn�Ճ�z���`�	�RE�x!a�N��Q�ۿ^�x���o��7 ;��"/<�#�
�W>e����q�s�h����l���I�L�t;�����-�x�Q�9��C�����qV�DϿ��kV{AVFw�}����F����5�6�na�m�;
=��f,#s����anù
Y�D�,�^����d�B/T3:���r�9���e};��)��a�4�����V��R��??��9ќ�K]�aGɬ|�N�GP��89"q�M@�8��3�B��}�����+��Bw���	4��w�4&p�{�Lސd��_�e��c�8�_C�LE�.WxF��r�sX���x�/�mt�dL6j�Jc�Z��H�4kw3�:��ǧ#ш��c������i1v�\�ORV
�E�H�����O;�n??��$���i�Y^g!����5Td{=Α��M��UJ֔�P����q	�<�	q��cN�/��1b�	�HMY�c�.y��S`XW�H@Y��m��XP�f[\�Qv�4�w�p�n9��3�	�=8���*���=�	ǇSo?�Ae�b�Hqp�!Y"�n�����v��a�d��qϻ�ISG�������������Kk��e���f%��Q߁�ԕ����r��n��� t-+��&��þ���#ya�Z�fz�%�7�S)�|�|�O@9��Cڻ�z�8wö���(�»0�?��G4���L���y���t��*�6�T��l��M���D�TF��|����l��.�eh�N�$��J��dW[9+����2sg��`��yo1�<G��	��S�ӡ)	���p@�����a�1T��9�"/n���v1n�g-���>��	��(����>��/9>q�긲\���eׅZ��N�4�'0���$�x>MK�kz�ӏQ�����R\G���PN�'�S?�9/����g��)�HD4��n�V,��V.?J��BǝX���MA��hy]s��l��"P����]�~���=��X�����j�t�����Xu��:��'�����H\B,;q�K,��	�������v��M��/��U&ٗ�x���RD~ݪw'���q^�s���u�>�Hコ��P�@��������.s�����uX`*.氵�M��O�'��e�H�p��0�)$G��V���'��1�o]�B�i���e� 4��]sP�[yUT�y������r��q�4�T�>ml##Y�-�Ó�̈���D��Iz�|��`����Y�nխU���r����E�l�ǳ�9Ƀ�US�C���$q�]�M�J��C�lZ�26}B��ή���=+�v������oq�I�Z�R˛z��W��;�ޑ���� ��n
��)��;�߰Cy�w_���Vh�����m~<}���7}�4�t"Um�8z���A�$�n?g��叟����Rm%�ߔ{�_o�!��4�VU���Z�_�߈ܒU��z���=�q�/�e���!_B�;��,�k�08��J��,�������ϲ��7e��U�/��e����w�}�O`���=���@5b��?|�����F�k,9�<�tk��HծnΊ��3�_�d�љ3��IH���
@H�Vl���
~2xk�0�<��ͭ+�e���s����\�H���j왇�~u�]�u��W��n�s�.������OFz���<����n_)�@��m��՝2�\��Ss��k/pt1��ī�R�Z���;}����E��9.��]FV��^T�֑X�
X���V�9.̷��{��E�@����S��-�����`����y����{x�͜��ۻ4b�m�\	ڠ�^�t�4%�[��6k�'0�-��~���e6������ME�!>�6������
�1�����cI�i�!nvܯ�#�V�O��W��ȅ?�oς����vJW�[��Wh����F+���9J�[4�׸�Up��4z^h���v���o/A�-�Y��/��~�i>�'
~�혃��K���9���E}9N1T�&�C �&��7��B.bpdHnkK�ڄG���caN���BfY�ؿ�&%;��Ƙ�g��w���;��Xʜg�o�_²hu��_�D>�Gh�����3�&��=����J�N�R��y�#�-�^my��6<X��3G�����G^q���v(�;.������p����`='^�=m���l���e�@���;2��ˁ��	����(>��򈙎3w[|}����&��*o��p��A[�5r�buE�q*_J`�W�0��g�ѯa�a�5�����-���Zâƭ.��.4^�/r�� ;��F�ia��u{ߣ1��	�������E:�Z��W��vr3�Z�Q�]��-;����~�2��\���!���Z,�[,�v�I����U�G0|0���jHY����9����s�m�_��8'R�&�ܰTV�/�fkl�u�:�ldX���vK�+r��>��3��+��6N:�0���֎�������ʗ�M��;�B{��o���
�}��F;p����LE�?P�������E��f���$3N+�6xR��9��֬��}���%ZҗBʒ�m�K�0��{X^�$g��,&�H�C����_��٭��a�� GVsT�wZ�������64�"��M��:΂)�ڟ�ݿm�hyl_����]t3)+����hⲅ����W{�{��_���d�>�ť���C��vX�ަ0�nTj���@�WF��x0����6�� �:ZIy7��d�5�[ϊ�� ��������U(_�.Y��dJ�dln���#���6�a��ʡ�h�Au��� �^�@�$ҳΑ��[��~�{Y���n�{�ƇY@@#�����8'�������	���3!��a��)qi{~-"M�T���$l��$frA]4�n%���}�Y ����!�g�5���(�����ˊ�{�o�-m6u���c>��G���^�{��^�[�"�+؀��v�a$D�"s 	@����K�ՏW�i�������,�7���T�~�Vo�~;�7�x'ԭ�uy�a�{u�����7`"6�ۜ8�VB'uK��N�2�\)i���*�m�"5�Om�=���H+�ݵ���@g����x��]ϖ5�"@bI�_wfy-{���	>+~G{�%�S�z"�����I�;����R��i����� �4�~������x4�"�<Wm)�tޛY������9ٖoIڝ�?�{�<���mmjvh�%������[����>�s�C�e^�mOKa˭VL�s�v$��h�Q{=�T�p"/][��ݢD�������RB�!$��ḒТ�ԙ�8�w`�����,oP注x���3�OS5h�M�;�f���5�,�G��TЋe���Z��.Dq�	�$�Lإ� �oU��� ��� v��Y��,�g�%�eٛ��%r����̮�� c��3�C$� Ȧ���y�ȓ���՚�F���7�ދC[�� J ����_C҉k�9J�a�?�߷�e�TJ�[��}�!�������uhwn���!+����o��z6|XNȞ�e$��hwީ`~��,�kb__E`_�����-Ɛ#hS��@��W�������35#�*�ҡ]�Y��cH����Շ覛s��>�t��R�T��t��\ìsi�.�}6G��ɤz�S��ᆛ�.l'�VWk���Rf���_2J�����&�H��%�����WM�:A��;a��_�K3���z�P�HT�p��\ܨ6���sڧ	���Z~���s�N9^ɀ�lQKod�\@(��t�,�9`�S��a��Pso��o-�t�Y�A�y��Bv�����N�4	x�4��~�s<������b��.]7�=kpmݷ�#/�V9^j�`�'o�]yn�.g��ī��e
��+�r)�c=Ք�C�eĳp�W/���'Vi�uxwtEU��?X�G�ܓG�.pF�9����������:��P|K�2ߺ��N_G��E��s��R�/«���lHC1��5l_s��Z��,��q��!B�{v~��&�,P��S��Xlq +�3��P�Ϛ�<uǋ�\&:*[�o��r���f��c<E���x�s���%k�>����r��X�`ren�������G��{Lp��r9!�a�d:�n���<�ܐZHsp֟%G/D Xנ�V$����H�k����`V"���_fw��!̸Y\�~OoP�G����{:G�f���f\�%|�q�z��l7[x{���u΁�u�y+	~{�oV�Ŏ�w
aK���Q�~�sγ��?M�}W����b�K�n�[��v�V��~�!�ώ�����Rr���%�eɚ)�����w&�����h^>��
yX9���nW,:gU��#�?�u��,��ߥ���br!�5���u�:ޥ�H��������[䲒W�	���nm����T~���������9�i�fLw�q8����6�X��VHg�����|��s;��W��i�d����x���r��K��0�d��YE~K�S�EYޘ>�.�[Ո]����{W"���SI��Hzv�F!4b	C�)����S)ڏ*�������H}�7�T��C���k�J	��ԧ���ŋ�(hޞ~29X��w�"�:˸��C��!���Oj�?l��� 1�.�����0t�9fحoj��Ҩ/�Yɴ�EPz^��xaYLV@���,�S�(v�͹P��>��u�G3�^��
���aB���h�f�3��b��?� ������/=�e����k��v���������w������+�"y��֥<cuk$�/�r������~V������~YAA{a�\岴���.��qO�2J�g+�q��7��;@�6��{�8Vp��OCGU�X�#	<��db�9nl
��BP�{�uNS���ɧ�g�[S�
nn�k5Z*a���0�9���q#|_����|�,�ȗ�\��C��Wy�XS��l4p(���ϡE��A�G�jD��@�'��S�,}|��&��eҁ���u������s���K�l��R�c0����Z%6:�"�e5�k���u��1{%��2&9��* q�tV�4,f��>��I��YǓ��_��*�N�m���Ut'8���x�:2����,#X�ZF��*�!@۳s.����#��y�)�q~Y�\.R	Kz�[J��J	����l/߭��7��M�q&�e�@�H�t;�}��e���s ��S���ڃT>�y����8o�6DBP��MV^%a��罼>Ԏ�H�>�ʷ/Ae��_�%/��>�1rh���-�<�%��ho+���L7�^���B�[
Z������*	w1�s='
�g���PYD��k4j��JHC���m?�b�Wnx�E��,ͱLZ8�L�%�Y5���n�0w0#�t���yQ.Q��!H�ѕ�L2V�I�(}�r��4�8����Lu�����v?��;��c���;���|&�铐@�0Y*�k��U�@�g�j<�J�Aa׵ 1g3��fvV%�FT�U���B����ZX�.q�IT����j9;B��0s���oB�RZ���Ul[��7��Rz���Y��r�O��W�$�,���  D��M�+y9���gdo��I�0˭�hU*=����F��h"���F�����БߜA#TI�]���&Ȅ�|t����L��js���ntCQ�E���õ����9�jʙ{q�t�ዹ� �a�$Zvŉ���,�5-gW�qЂ�
Ĉ#�;����}���*��P��Ov�[Dım�����6�z�m�&wH�ݩ�nS�����ۏҁ�'N2�nå�N�iy-cҗ�����|�#��Y����V��HG�ִ��A�!:ɀ��n0q�/����z=�l��թ\����|�)J���O�D��sx堙�Q�e���[����F,ca�5��a����l��C�ÉV=��b&�ӀQ7f������@�:3���c�̘>���=T��vZ� @7��ѷ���o�|	���eO�}ˇ�tm�D�L�rZ����:FV?�v�KP�^w��u�#ޡ�G�c�>��[H��}k�O���� ��f]d��]"e���&�~\n�q���C��4b�XN�|K��(u����_9�����|��Nn����!7�;��+��<a�l]{�{�{A�'��[A��P���
3�X���t8��&w�=�[���gr�#X���>�Zn���X��Kl����З`�vB�ĥp=G����GW] .�eP���(]ĵ.f�F����'�LF��hMGK������ݠt�mz�5�ض��*��Ѵ�(�g�ȸ��|���r]n���!<�Vq��m������K�� .cN{h�����o���%�9�3�$y�9��S��f�f1�Z�%���qb|�o#�'T�#<X���IG��|�a��Cꪔ-�rW�ʗq�WV%�N�mV����vx�A�����B.t�8�<Bs Jb5�H~��C_�q\t�(�~{X��}h[�}*2{��+_tu�r��B�����,i�-:U�<�S��g��$=��ß��j��ͮ�nR8T��#{�m��lƛX�X�4K�ړ�*zo���p��s�lC��ݲ�\��a�us�Vtr�A�_&sT�?��[�{gM�`��}r�����%I�j��1zo�����Wr��9ƅ>
JHi�&��/|����	��\����X�\���V��2{}��s�>�����=P.�1al��\�At��$���b^����]�٦��-^�'އ.ZyK�Lt?��8�C-�_o�`7#�w}��>�yeE��������nW��~N�$Ip�<f��	Wm/��՞���K�'2���{��ޡl-���뵱.݂�V�.��`���>�Z�g�_)�� T�(MT�;����wv�����{����@	l�lp4(���:�%�����c���<&��,��Q�?0|�Ƿٸ�����s	$����].Os@��e�����1�l�JL��vkg0�d(˷���*;�	x���7`0Y%���Q������b�U&�a�Ж=e̟��O�����^s
]9�����~H�$N��o�YQ�o=P�Br�e����E�&�C"8T�HZjU��`���ͼ=��=X=��A��PTI�5�#n�Em���7�9��0�(+�Y�D����,�Z�&"7�iΞ ��Fg�Z����m���
}�[q�!"m`jA��Y5�_�r�Mz�u��\��ѵ�l�Ar&c��U������	���x��+��¯�߁x��d!!d*:�R��%z�75�O�{����K�+��=�5��0'1D�?�U���S5z[b��f.É�6!�ニ����'��I��Ŀ�h��ŧop/�aKl���"�[��V�J��Sz�FJ|������A�����v��@	�u D���[������5i�������ު��r5��VۍtŠ�X��}.�����6�>��-l��%Y�tܴ����j^���yM ���Сk�6ǰf�� g��JL����{z����h��L;q��̹\���cE��r���}�rw]�X7g�P��)��*��3���)J��Ċ��nz����'��5�h��G����ҳ��ے�\�R`�~ш�M��0rd��C3*}�r%�O8���9�o]��?>���z�2`��
Jǌ|��ȳ
Jފ��A97�g�^����rs5_.�^P�ҧ�~	������?R�O��[:Gәk��p
)j�0{�ȓS��;�g���W
�ȅ��X:�ZV�EI����sܮ�K�D/b�^�p�(h�1�Es}�f��zV%ċ>St���r�|��߷k�[��v4"����'��������Y���*bȡv��-Z��Ӟڨ��[�������j5���Z�:x4�(A�Y�
S��gn��Tճ�8����'��63�r�]t��h���Y;l��?-g|s��M�H7�z�g���tt�Hh^u�
1`����'��,�TᎭ����B��n�U�k������l�_� �쮑��Gx�1
���w"Py��ݱp=�j���� �|��f@ƓſP�k.2\�)�"����6��9�?����	!�))�¡�ݦ��n��h�	�Y�T?�XL:x��"W�-&#_��P%zs.�0$1ƵEx~!ベ4_��k�J��C��n�*� �?ȏ�uH�E��u�v�#G"��0e��9�؅�ˉ����"�9*��q�7��{5�s��r\c�����X��+��bj���)��F�r�E)%U��[�<v%d9�}��Gu��M�2���4�EN�����1�m�#*������5�h`�Q��[Nկ,���7I��6�):�4v���'�o��
�t��[�..Vʫ�����1�d|�{����㉰��t�{M��D}��\I�S8�X�1�?��q�ݱ�v
\���3��Ec��ޛ#NR<�o��D�Rf��Ν������^ �� X�L̯m2��ـΞ
1X�p���M�l@�{�U��M�]֠�W��Fa���?��7Du|a�z�Z���%�cK�ө�>�������~d`&��k��o�g�Fй�`伜"~�q|fPWPR�%�/8*��Y-Ud�t�JA�LN^��U�+��?Ą;�>�X���f�������TǥD��'̼�:t���f���=�o�y ���Ӯ?�x��5�M����]�+�<n4$�Cg}�#$/�2��o|`!�\?�nvh�v*(H������ejKi�hx���d -i�.,C��R���l(�b���v "�7��W@*��F�J��Z��}ώ��jta��	���C��yB�����s��G/�g���5�m��2�k��w>��D��1ս�����_�g��C��%l$�kj����m��ɳ�y�����w8����U%�{jj�M�J@2�H}S��{��ru+��?���ʶ�D�NԡUZ�&B6����\b>�H������V���D7�����5ȃ�����/��I���s"�z��A���6T~��U�)�<���׀�ko��'���Y�����B'��}���>4��y}4������ժ�T\��m.�<���LF d�Jg����@��]�Y��]�	����C\���!ߺ7�Ϊ���}� ����P>�Pi�s���W21�%�Jv�x�JJ�=nm���2+��b���%�b��A��.�Ђ]қ��=�-�YM���j� �D�څ����B?sŒWd Ƴ��|���g�v�;[�ye�l��q���h�rf�Î�C�V��5Xt��1р��;Y�� %v"f/��pα��=��[�[�ia/<�I|��YPEvy<�T����%�4S�4�&f�4���5X�'@��*�����"9��Jf��"�BEzy�[�-I��y��� �4Τc3Vw���UӶ2��:B���6���w2ueLH��pEl㽽���A���,�,�rL�8 ٔx�T9g�+�j�S	p�oA2��L&81�A�hP霄�U����]� ��#*�H��5N�k����ÕG�8
�N�8�[�����}j��W��a��B�w��t�̽���ef�w���	�~��!`�)��WA���;
����~�w��6+�^j��0�-J��3��SC�� H��R���r:���).�?�ﭩ���}4�Q]�W�K��YGM�$ZeQ8�"_R���1�H4���&�1��s��;���k4��ѫ��QǢrG](�-���zIt�J�Bp��r��m�r�A0�0��
��Rc�Y�B�<�u����j�{t0%򪳎�Z�k��$f%Yc2<�l'|����{N+���3��ԭpHv$d����d��Y�cv�-B1�W�a�6���ND���N�+���n؝s�߈u���A��&��~^`��P]��k�r�`�J���i�SN����iw�s�T����(ڪ���_ݤ�w�4ɍ�������En-���m�sd��c�ç�P�g�2�:y�-,p{U�t�%�a�#��:����L@��.�+���`��mƺ�����[�(�T���"�y�����_�^�%{!n�}��s�����ǡ>[Z�I
/g�!�R������efA��}K�ב=�K+��}�{�r��[/o�ՙ�|y��?<h\��=������`j�A��C0kd����NS��X�k����߬�[#�R�+��a�|��p��;��A?�'��J|o\Z!����;Z����������J�QX��i�n��j��$�����?ͪ�~�>/_�T���J�9P��-ҍ��S�N�m�?8����;�N@Q�j�x[�N�.���͜��#:~J�� �($i^����`9�6�9K|���&��g�^m�`6�5��e���fN��ޟj$rsL3�N��M��F7�*w �jVN�#'~�T��X�,g��t�K�*�p\S��f���j�������H��ﷸ�@����I�A<����(d<�b�����L ���O��l�Z�}��[�h�5i���U�D�T!�L^,)\��,�?�m/d��ǃ2�u��jʽP��Ԑ�d_��4q�ȡ���u�Z��[X���I��DD�YW�@�Y��Ѹ�{,sa���6]1W�<,Cr��~4��ES����bE��Ep<^�^=��|�I�LL@�{r�c��q�>�vm{y���ug�ƌI�gX���3�=�(��A��,7���͋������L���#�e<��8�`>Y�,��)Y�5�6Td�pV�Z狳��~:^�	��*[_�l¦x,��=�|V{��۠�X�}�n�F��W0w(��A�;�U-�v���s6�D������kA)Ń��$����b�Y���٤�T6w�`L��^��}��⼙���A��2~'�q�����f{���}K�����~{g2��������{��-̅�B| cs��'5����a]�XAr��P� �ڷ�d��BI{[��ռ�s'��~�U^z(	�7!L�{�eOdڭ����������kwx<p�C��Jz$PrdE$=�)�t��s�o�[��}2/�	�=�"C)B0�ȗ��\0�OT�Ө̩��v\(Bfgs��h��]w��~j��7̶���w�;�)�pl�F!��F'��t�a֠�?Q�'��	� ��%E��`z���>�X�I�*/C�٬dyZ`am
�?�\iUp?�O�qc?��Mu�p�rN����v�/ó��ݼ���)k����wX-\��BǗ�m�y����PFϿ~t�x!�`Btn)�U�﹐�#�v4��y�Q���<�&���W�m��W��3�NJ���U߽{��ks��{;�ҳ��c^ GҮ��`����T�rR9V"t�#���L�T��}�+���|܈D\A�2�{aq�쩎3/
aB��DBZh_��Xо-'��m�L�oފ��w�� ���Ʃn��Ko ��f#p���5 H�2��F+�_тu�dV	 .�q�.I�$�TqS��E��q��,;��P=�Nk̻?�2����ݣ��쏛��<��.����� �?�B�)���-�N�7�f����R7�m��D`����,���u}�]՞H�Y�U^T<{��EaN$���ƪ¯������nU�aq��.���`�af^7��cڔY���1�\e!e|�%���@N����?#4=�b�J�h&[��J+
 ������z�rf��	*����j!	�G�̼�ᣉQ�y[}VM�[���ϒ7b��DhG�%V�E�ۙ�.��!�=̚�=�	���æ�5��l�K�����&\1�O�N��Ժ=�Q�|l����/`2��t-g�)^��yW� �LN���6�)RS��㫪;R�^Bh�l�E�4Φ5�ƾ���x���f�]H�ٖ(��$��m�9�7��^(�n��ܻW��Eg/��ntpxA{����e��5�=���Ͻ{���G&d\jIȉ��Sq�*;Q�zQXߋ�����c4��L��N���:�^����1e����W`%+�C�q>:���)~�)�Ѓ��.6��^-�uG�z���[rdJ��������4���(����|�E�}������G4c ��jO��ڬ/2(�f�z�9��y�ި�G8k<@ȖH��Ԅ���W��Ng9�Fn?K{�����q�0zmє���>w��m,2�g2C�=�i�;'乹�ݕcm(��zQ嚛Ĩk�]�ɦzc�A-�x�LXE0�L�Q\ ��=�$f��]��K#�qkҦr�D8֕v�����rl�}|������^�}�
~�����q'�"�7�
j�:�n�ۜ��-t�<��M��h�P�S[
�xN����ns��aV��Kٽg��W1�73�ZP��GA��+�*����[�����|͡�6|e}��2Ѣs|��Yj����>���B\��fA �؞���T�u$r����1 K���vY��m�{������<;d>t�:���#�<�M���Y���خ0���F�;;/���g�
7��	Z\��!���� �w�����Җ�O:r�K���ũ�	����Y�,o�G�9\�u�\���`���1x>����u���oʏ���s�,��Bl�J�_pu��=�!Y��j�������@g���?���:��������G�D$yY�oɋ�n�j-�okR����ۉ{��ҎL�b�(�?]x���T;�f/�{x%�u��`<T�ymcV�սZ�q#�/�ƙ����'<�p��N�C���=WexP[�H¾�sy J]�tߎ��m�IL�6r�o��#�.`��w�������=v`g0"�X����V7�޻6�j[��=�"#�}��i�E�ŚDnqA��
_z<t:�@*ͱ��`���q%m_tcE�U�s^�í�-�^��yq5
��/�#��#����H�fq-���#�7$P��e,������b�,ָG�Yc�GD���J��G���=}�W$�f��(cw������	��6����,��H����h�i�֦Po�[u�V��"�,�e!�T��8�x��_��u�n�po爠�r�	;�����{��?愎�����-�䰴ָ�螴0n��E�����K�۬+L �8z��6���<8s@ͷ����Y�;��{�-L
ⶏ5�T�#�	�KbΒ�p3�4H�&S��!g������%WTB�#�29읦�����P%!���\��5���ݸ��j���V��i�?�뿕܍��P�
C *�rWr腸)���8�x��wp8�\�ܖ�냪з<2˳�� Csl�DJ��>�B|�^#l�+Au�}����\�[�Z��yj�Ϸ~����������8�P8��˲'�8�)����8���c���Յ�Ktˬyxԛ3�!w���E՛�ַ�|O(>
�'��!���1V�!tt�,���Z����>����^��2EV1F��1�}�T���6BT��n���|���j���^�J��Ժ��P�B�|��{0vL���)�:2N%��#1������&��?j.�1
`�^rgZܭ�+��L[7��S����O���`. ��pVP�[��q5�D�Y��gM���|c����v����^�~��'NA� ���~��L����̮&�Z����@/0�g��4��>��>@�[}�˩�+d��xm	dK�,t��k�����}�wx;�_��r�W��Ug��}t�	�Y�a�e���(差˟gC6ѳ���A}�,f�d)C�Uҡ 毖�t[�hb^q�x>��._iN$��\N<���r�,�,*kb{��/�a,��]���Q�T'�nw��h��'<�W9ָ���D�����>r�6čJHe��w���������� "�/�2��$`sXGq���׳�7�6Ĉ����:8_@t��WuΜ�ω��m�u+i^�`��K%��he��E.2�ƫ�*��.}2R���8�r��k�8��F��ȯ���fU��6���j���_I�Bws[TOq@Y�o��U���!j�͑&��7Xk��F�9
�)�v$�f(p��Ob.Owk���%��nю�6r�t
e�SzU�Տ8�㑭�h(�"UpQκ��:G�9��-s5g�����p�ۓ��pKr-h������d�T����2�WM�O7���|�+�TZҷNY��b�� ��������u���b�ŋ��"���ڷ7��?�9V��\�WR�Q���
��C�;���z{(��{����WZtV)ч�{5���4�/�����iI&�#c����H�<�o����jpp� �̹v��Ȅ�,�ù�;��%��B��ő�����w�*l[L@4n��{�e����vߚ���#`|K��n�$����9�Y��M�|0R_lZI:�)�Z]6���
��[͉��#�g��h���N��`�&����{u��v]��c�# ^�$�J�ps��H��-+�l��s�]�[
Xϊs�Y�D��J��P��+#?x���X` <���+F�W���n}l[h�c�߄����/L���n)V�۠���t���ri�0����>�D}(U��pQ�V��v����a�����Pr~5���<ݴ��eFRҫ��^����9K����1#�IFe�-sn�\�m(N���.����ct�`�tl�Rܭl����d߉�GY�? �#R�2���M6�qUas��x�V��+���,/2R�P+���l�� �G�����x!_��g{M��؁�fA�,��"[WY���������@.�ڡ�	`�F���h��=27'���m��?�c����d�f��a���T<���~���mχsH�!Vx�⨉��l|]��G���HF��NY�xl�%wX��vʁ���	f��~�ly��HU��u�3���T
��z�x����Y3^7�N>g�tZ9)���S
��x�j����}���^���R�~�AP�X9[��cVM$�?s8�^��J��͕
lIvs$C;o)D���ʸ1��q],T�
��l�\��N�1��w��/-"�ɲA���@���/aOB�ޡW]6TG�=3I��8ҬM���JE�"Z���.���d��
EK^��b�c��6���r���n�C�(��H[��g�9M�M��]�`6{�x�&Z�B���MS�QM����ٳ���'nְ��O���5�m�����M܂]A�+�:$�]�7p�N��=�Ua�eL@��\ϙ?;�R���T�s�hD��%}�G�*�%v�����%*�l�.�ż,螝>'�OF�����$�j�¢q�kq�#�1���'��hF?�8Z��y�3��GU@��j�-v���ߙr�GC_9�b��Vӱ� o2�5a@fy��s;͂�WY%|��즫<
,�5�8l�J���GQg�5���<����=���DLE���������>G�?^c�,�csY uN�5*y1�/ ��(tE2/�7���.��A���k���):�ŅpS7mDCj��
>��9㼅�+~���?4	--3�PsS�]KFV�մR�>:�J`�$�xYI+Ԑr|r���[M�����t�6z���Y����h:o��^����`��R�9���"��i�����3�IE����"�X��X�-��ΓD�EvSr�����f�������uZ���N�w |x����
/:��1�}�+
�]#ٵ\D���2�6�"�,�2ke�ZxQ�:g�\o�:U6��Z`x��� ��9�䝷��A�oo�����U;b��mC;��sH~�_%[�7����T��w��n�'��] ��҆{��T�XIK�l��@���7ا���+�Ӎ?�?��O��x/Z�����~㸷#}֜5'�����GE7�{C���r����v�s��)B��Q��i�Y+��?B�>i	�(:�g�����
ܝ�� 4�D��]�H~7q>!��}�?ʨ�~�@#Y�b�Nؠ�.H���G�����Y���!ƣ �U��
����*���շ�yz�B����^���W̆.������fK��'2��\o�lN���\��ek`ao�`]��Ԣ��
�#Y�^�l�E��X7�\$n����&�7��f+'o���>%�އ��Yg��w3�%b�1IX���_)����	/a��Si��x���|Ѓ�v�S/��
@Sތ�{6ąP��v��80*1:5�y~����m&��xm��q��87��Z�/aV��vN"���i�/�x[ ��b�t%Ӹ.���">��
���$���P�S{}��x�8\z���'I�{���/�uv�"zO�9S����#���m]�i�|����뿍�����t��$�n���j���5@V�<�Yݽ����IXY�	�{[v��B-N�|ha}nW���xC�;��"��\,n�H���'�8���;(g
6�+[���^X/sn/.O��@Nq��S���zQ4�J!	H@�|���	�6߂�}3���B��&
iu`��	��+
O]W�s�wa�)��F��ۯ��c�4���M˶Ic����&�e�I��e�#j�+�e�,%���(f1�T����K�B���o�.�j�Ttn�ִ�A��5��B�(0u�0Su~5�[�TBP��q�{���v�0_�2��^�[��yA������'�X�h׾�/����:��ܻ�L�;@=�:'��9�T��ݒ�NnT�$�D�P���,��o�����j�m,o�(1����-�dF��s�6��=U���5��2����e0�-"B6	�_Jy������c���^�������lU�
ǌf�TxvP�bk��7R�a핁��̛H%~�����Eo:��P�Y�@����h�Η�����e�w'��8e��z�G���9�8�:G	\q���4��Y;soφH��q�::��"��?����Lݴ#����Bز�=�c�`�fa�W��9&��5�j��-�.nۦ��)��/cdNYC6���m#}n�'w��]T�q���'N�F8��z=�������?r��(6o����t+�D-"wh��Q��W{@;�o�O\�bыӪ�R��%2�.a)���"�S���M
�5��8D�&s%�B�i}p=���J�߀��Q�o��x��fhGT�@�WD�t�!�^�)�-폈�^@M�du�z�	�yƮ?������������
<�@��?dA�OQ[�<�it�L$>�����H��ti��s����e��\�mR0�@��(ۧ�a���;-�������eE��#�bYH3'����?s۟���=��Z��Y�HǦ�%���P����Jt���'��g��'���ݒ�A'W%�5H,n�Kb��=����f��#z����v��9k�z#��� ���C��
��7�ǧ>����%Q���������-;@�P��Ȫ�9eXT�9��J`^�e$�P�6W�R
��7S�я6�����*�4N~������O������I�!�t�p]9j��:~/e�ā�ǢO��{���������$��lB��d&K��s=Q��or������'e\��C��$ ����Q�G���W/�:1~۱X���mU�Yd��<[�;kVo��L2���9�O���*m�w�S$���0"'ɍ1��U~�cģ�����YW���p�IJK�[5�ƾi�����	�8��@lp���"O�Ǭ��x�֤�Nw�FDM����\��T�s2�/�*��{��4ݲO�~��C�7����.�J2��8�{Ţ����H]A�[!x:���ǳH_?X0�<�%�	}� hI�)۶�W@\��o�?Pe/���ԍ�"�u'�;�5|P���s������"�%�V��$��}�o)�0O(Y������Q�����"]6X�F<q�V*\ڷ��N�[m�Z!|�f�CW��-�^KR��|۔G��kL�W���2��S]+�����F�
��c���f��Nv��
��N���:�o?|_zt��A��!��moHl��M� �MUș��o$\��{(��Q������Qӥeʅ�jkS'Pc���MA~����}���_�z/����q�c� ���
_!��#�����5�;���D���S�c'N��f/�	���y����ț�h�jH|QM�HO���W%QV��W��Ӱ�qB�*���VV=D8mD�`�x�4��"O���^�b�U�n+�T֥�I�1�jb�-�H�Y+�/��߹�q<���EB���a����,��,8D���&��3�����)la��.�zi������f)4�\x������%���h�����@a���n�tx�ϗX�� �9ՏH򲟽A�b��'&v�'4����Y[)�S���Ϊ�)'@�?�l�C���<n�n���'b�>�קy��0��+�*��të�+P����z�2�=��7�9�߰����e]K.6&�p'��+���˅;�~?����qsƈ�R��o�KOͷ�z�f1�U}���H���!��t��*A��ċ����՜����J�	��(,��m��K����=5�A�� u;á�(c0�\˽�ru}Fk=���)-�[���K�������k��^�����a����ā�;���!��Q��챫��V����O��5�E���Kڱ�v���@���P�?2�� [v=L����G�u�$ɨXF�#a�3O�Ϫ9k;�jW��
��0��X�*�����6��qV?�JE��w=I�_V;�7N(�72 �-�b����B ����i��\�X꼗�M�dP���g�9=��/6�7ϺA�l�«4���y��PS����|��z�Z�s�� ��v�����,.ɏ(�;���\�	!Нy^��W�'�𼹁F^\���ۯ��C������ܳT�������IJ��j���a���q8�r�hދ[�ʳ
���HNR��ܾǙ���qy��뾽A��Y��[W����>6a^П�z�^�){@PwSڻ]��>���Ô�'��Wa�P~��՜����%#[�:�Ӛ����s����@���o_�S`�=Ջ��(��	��&j5Y��.,�xN����{}'L{d�Bj\��ü/xEM
��l6�Z��j�l�u���kVߢ��l֟܀:Jʬ\� @��3�y��GB����'ƘB1�%R�{EW\ȗ��߆Y=��ͩ������S(mAT'?7�	n�����tS�6�!EO�5DBz3�P��S�Ok֐Vnú�9E�I,\����$:��
8�bM�9橵��?��)�{Q�%<u��Y�M<9o �I���ϯqYYUzr�F<4<S5˶:����b[���z~u�C��L^,iì��%���d����<��j~���!��eJ�������	��G*���x�.*�����Ki�Mr=�(6���¹8�@�_�����2�"��' ��������,��K@�x�89X�Y�U�6�P�D��Ğg�bVc�@߳�Ҍ%�v^!���[�	J���&�ߣ<���;�{:��ƣW�g�Tm/��;mk������Q������83.Ȓ-�, $�RK<��$�/��F�C�������p�G�P�J�Uqk�LТR��7�G����$�2A#�``�ɥUmT��W�M�d�W�j�|Q��.�i���� ܭ@ޑ�v|:��jVv�WB���^����q�d��b�=4����%/�������&V�x�*�tV�V��h�9>q�6�X���|�En��3�dsP�d�֓v��x�M5�+m�,7Xח���@�*2HVD��;!t����x���p�b]�Yw|iֶ�Oh�x�7��IɌX<a�D��v�h�;
s���}���A��DI^�*�Z<�r���ѓ�}�Ʈ+��9����mOɃ}��h@�W�r����]��01�h����~��]�=h1�����rl�V��s��uQD͊S�5ա��oQ���pH���p?����������%�����#��.�(�d�"�`G�,K[I]�ԭ]�M:�@���6�'f!�-D6	�l�h��%�G�g����+���5�LG�����|r�T<���0'����RN�:��*/�,�{��EĆ$�]�1xH���9�����=��jX��}�&���'4���Tp/kv���A�hӮWa��b���*3�o�)R��i��;c-z1(*��ص*`@���@��0��h=<K��8����B�bQ� �zg��m���
���?������h���Y�Z���
�'V�6݄�J%>L�M�w�S8�zY��[�Ԣ$��x����7�������G�����q	��z�rѱ=j���D������F�q)j��<�g-��xr%�F�l�:��sr�w���3my�&�%���-[g/��mr������C4���m0����[�`؜� �,Bq�nΝ=[�������羢��ɢ`8���.�� ���snͦX��$���0*b�+�Kk[o.��j!@�fmS'�x�ԕ�z�m3�̞hxE�5��~�%~h����>��6!VQ��2W�%��0!CvS���Y��縮���V�|�ō��9���ϻ˕������Flcx�M%[�%}�,�rN��xE�^���!U�C1l�A��Ek��B{΋�y��{<M)�����=�wR��E�Ű�e�_'�����ݧ��Y����D�{�ֈ����m�9��g����>ؘ_�uG,��|ݑ��T�Z*��9M�p?�גK���%����,�6�J��+�x!�/qOTM�V��K�\F�#e!,��p4��3�I�������Ja�^����d`��b�z�j�n� �=��Mi�l�c%)w�0�F'��w�|ͽ]��
</(��F;/m/k#�ꦸ��Q�Xݫ�yݠYl��w� t\W�T�G��5�1=���r�cx��WzZe�*�/R:�0��-�b�eK�ܭ}c�0�55������ߗdǇ�%JqQ�i����!�u���(}����/3���x��4�8l��Rš|�tg�������풠š��
�>+��ꀧC�o�	���{t��Pj���tPUގ�5��+��^���\=���Wу���p-$D�����agg�j�z'@��hNd~���"���^ Q��ۥ�ܰZb��!ޔ�������'1�
ʷ�O�MR4��� E6��/Ә������)-
��%�4,e.W��7=�<����=���T4��L�>�j�%�Z#�;�0UUT�E�Ƌ�Nv����v��7��)�]���1���X�)�Y�"��ER�Y�ɻ'��9��آ�DꏍO���	������-���)X?Ǩ�u��a�G�kTNY��'+5���豜�D;���V���\z|!������ ^ul$�3BnH��ss�X��b~�J���I}�O^��F��hVέj}�X��S��/��`�o#���q9��mhuiX��*�@�'�f='����Il�ލq�`���N�^��|��7����������K,����+;�h �=����r!>����Д|�� ��>�6�.u��
�Ŭ����x���1�57P�
pC_�5ø���7����:���q�=�fh���z7HL��yTV��5q(N5�Dv ����rkbH�s0Ch�#fL��&Z*�T"o��nťi��r�@%|�����2���6������hD��b��?L��Q�+zH��[1gl]�d��֚0E���n�c��b����]G8:?b�	&���fqJ�pT�W!��i�P�<�i��v���zJO�!����q{ï�Qɋ#�����Z��v2����6��,1yL����:�*&J�~��}���F�^�lh|._��7��}/ ��^�j�����g��͛������]࠱ 1q�ҫ�t��W�6K^�O���ON�{�:kܺR�u�ٷ|�v���L�QƱ�OQ�q��`��S*�C�2-d�!�7��Ē ���Os�oL�T�T����KI�E���:���f�oclD�P���.3�O`A"�-��gjB��ޠ�Eތ�p��
��uJ5#�!2������:�: �;n���Big��5�I��v�;����ak��Dȫk���e�)��Ϸ]�w>�7����K~gFU\�S�׶[��� �"�S�m��������~�/2d`��0f%pr+�t�/�xt��3q6�}���"4�i(,7����.����^)☝:P7HI2���J�A�ì�����Z�W�3�J(] 0��s���&�e�w��,��K��Nq�ȉ����
4 -��푻;�
�c��!��o5�k���9�W4Y;r��W����q5�������0��'�g�xoj�Y�;q�F�y��N���)
鱵�)𔲑��(�mw"ݐ=}+�b�͛�����g�,���I�#�]�~PZ��8՚������}���G~5����
G���a����7k��c 7�G��5��+-�8K�欘�19t;��Q�:K�/���'��K�	��9�=�V�`UX
�����&ʣk�Է�Z4��س�l}��+�� |�lI��Y�vS�����{��g�њ��!QE��3~s��� i7������K�j�\iI*���j���w�i�_��ÁM(O��� W�;a�
I$v�MM�=��P�?)|h�F'���ix��v��82R�Hr|���mХ����9#�{���a>~�>�t�q�:.;�z��\W�56�Zt��(����t���jB)�F�Z�nZ9�tߓu�l�3���h��Ʀ9�'��w��7<&��%"�'����0�Bc�/��,1֬�4Fz	��io������W�>��W��O���e�i+�!����K�9H��`S<B?Ǣ��/w��u���j��*�oZ&Z�B�?�?6��"x��S�O�����w��
je��q]�єŤ�jN����xo'�9��B�-/�v�i���ΐMmG�X���jh���c6-�n�u� +�2o�]���qwH���1t���O�ă�-h�PRs��v�r)��9狽b�y�`�K�|��[= �Y�p&Y�J�8VI8���3ߓ��������F�����M$v|F�����Ւ�>��/gQ�;8=�f�k-P�"��Y$pO����O��|��u��>JX�{p��A��`6E��2����ȩ؊+�ƩF�����M����i������m4�YV��|��g��K��p���z"o;pԽ�x�>��1�w�V���5�ʢBb�h��&��+��÷q/|�ڕ��J����F����F�����/��uu�D�a5tT}8�b��m����}ư���_��U{T�VN,��x���ś?d9\�{��m����U��_w�Cx;�!O �%#�|���̿�+����W �=R	������3�,l�e��۔��2�߾�?���'X/j�s��Y�qˤG/���6�|H��o��}���h:m�CO�$���Sit+æ��%X�Za}��|�]),Q��h� �{N��Zտ)���_��
�]iIM��6�o>�6��t�Ϲ4Y9o������*���|��{M�c���Eg$��|\�_>�����u:����Ð�	ku�����OC���?����N�3|��G��oQ�ė�8�r���sN��	{���s�����W�~u�vO��e�p��m�E�;+gxN��ܟ�=��W�3���I4p�����h�kl�i�w��ى��#&2�?o��O~��봁���nS5��.�� �ӎŮ/̜勤�:|��ű�r�����rZ��Fڕ����Y���]��-Dfis}ÓCGS��P��~k�?�t�{O���s���.�[�Z�ɮ��9��>��ǟ<DO�|���K����e:$Z+�m��et5�׎x�� ���#�oc���do����r�S����S%u��H��d�����L�_�������>�h��q �(�8�\��</_��%+I�mv�i�����@{+�ڣ��)ݏRQ��t&o(�{���,;[��n���%�9E�ϭ��ηۧ�+gh�jp��v�U��9�����R1�sW���t�3���v�9���X�S��1֤���}�a|F����*�;׼�Ļ�re�ʁ�T|�(����O��W]��r�w���-�vǪ���݁��æR���ٺg֢���Y��*��rfI[|�������,��f�*�O2�&L������`�~�K�(�pi;kA(�#��}�_.�%�]�v�K�{Kj�q���BӼ��8p�H�)�|��"!�uO�5�ߘ	_���Tr��v�V��p��km�/��x���ZJPՆ�g�p���6W{P��ژSJ�c�����Mo�u��H�~i�ֺ��ZGSc�w����|����v�hc��Bf���2&5���bV����z~񙷼��m�B!�q�Z�j���h��	��8�o�����F�6�M/, �f�O#�̶Q���,قo�$��nB�,R�eEH�:[e�����h��x�W�P�x�G
��.��%Ǟ;5��|b�?�&	}�8�ʊY��#}S՛�l�ԩh;�7�@X�i�b h?�1�t ���ڏz<�����%���s� #i�K�M�.��Cr���,�����^��+�l��bN����e'AA^���m��8L��!�0�t�(M�ݥض�y�3v&K�����$�O��-�����9��9��Nkӿ*@���+��Un��OpGC���	,'��3c����O��s�0Ɋ���Q�rG^���b�:����y<Rl����i�8�9+7u���8��E��B�?��E��ƀ�z��6��P�VD��ǝ\�v�����Z&�y�����<_�8T��<�O'�F3#k�Ѳ��[y�a�Y��������,�/[x�i$�tXβ�gC�ޯ���r8(�pur�X�������Ȁ���pR�EyBk!;�7����ﶙz����༩�}\wW�|�n�Ǻ�Fh�YV'%Cދ�(l�cS�MKG	�<;e�@�ّ�؞�M�X�x�ڟŅ��y���*�Φ��/3��\�PEo��?��	��ZZoSX��� ò�$�9��{��^)<xW�l�ވ�G�����t`3�=��W���Ind��g�9,p���na,/Cq!���V�仈�:s�k�q�bf��#��,��Ac/@1�30�%�syoB�!�nl?,|�8���v8�@)z����'�{�f�9츛��� �RB*������ᚢP�0�/(�e@;�V�|o�X�dUe��y0�D����Ĉ��g5�'��8%
ɵ����X�/� ��y��݂`�*�6,�d�$���1ǱpX�W���'V�ՖR�:	�}�!��MQ��*��H)wC��[7u���<��X�uKO��6K��5��K��������>���c��GYdX��*�d)���XK5�)$j��cC�o���� %0^b@�1r}!�u$�`��"֞#�O����a�[�_8k�`��Gk1�@��f1M|��j�}�ɍ�c�ج(l}*�y�*��8jVg`Zy���pE#[�k�n]\��%��4=�P��q�ӖR���Z�\D��^o��/�� �ů��O��BY\�E@* -_im��Bn��1���x�4��B�M�J1���E�Ex��@���$Y���)�ɞ���^_Z��U�R"٥sZ��`��\<�M��7�f������"b���RvZ�r��k�m��1	}����)�d,�Pd*��J($T)n�4(���G���%1��:s��\�W֡���'���z��S*�KY>!��pI[Cڒ�ز���U�5����9��6�{
�v�;Ӊ�2$��{�Y�μ}����o��q'E�xto���O���k��HS��b�U&Ց�hv޵�P;�^��]�9O��s��(�t�66�@�J�%��)�ռN��տ�:������+��b�� ��MA�&�?�gz�|D�ኰ���A����
0F�n��b�Y�;uS9�+Zv��e`{�)���N�PP<ݡ�~������{ 󧆖]S2�Nڬg N��A���9��J4��A��0~�7,�u^�:F��1��vS��3�H�^0���EDT*u��+�;|�_vs
�W�����MA��Jj��-�\�~�����ƛ���}qOmCzh�"o��Dt!m��Q�����4�t�~�澸(�����桂����Y�y�*��v��p�s�b� P����Ԏ�Z^E��N�Y5��*������Å���~��!�<��
bV�=.l�ޗy��̳fD��������uc�~�8wSK���O=�x�خ|�RB�kn��{`5￞�{J�v