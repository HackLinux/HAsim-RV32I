�ƌ��TP�f�t4�������F[�a e����@�7�'���pa�]�~4A��kB��I=
.��"O]d f�<��� #0�E�lJ8��ހ�5� l}�Xj�����&#�x�H�Mxf�� ��}���7�`�j�FK0��m��k��~���En�eLr�	��~e�m�@ҿ־����1�J���!D��E��A�4�s�%�����0d����
�<�>B�D��I�E*?xM?T��3�q���c"�1<xB��Cy��P�-�V����}?�[L;(�a �XΟHlYe,�-��V���:�c��Q��G'n��{u�r)d(��V��#�`%��K� ��t��&�J;���݌�'\�/��	���2��?��@��g�lL���a<��Ii,ST�,J��d�@HY�f�o-j��k�K=�Aye���qjҊ�+��O|x��-����0�i4�k.S>�tk�)���UBE`F��R$\K}k��%����w�53�F���<�Z���i{K�=��r��pn��dsQ��J ��M�R'?ߙ�
�r �n�������fj���B����BK�6�VX�f�K�u��)��&:9	za�;��]V~~9�v���CҀ?;�w�7�e{����?��`-W�RC>��^@���{��缔��uo�H뵢�V�x�jE���s��� ��)xØd&�v�(T�>�����At������2i@�@䓜{�����|�e����hQ@��_Ʃ�D��<b��f�VA�p���j��L��� n�l� ��W ��V����yb1xg�J���{��p	�P(�2���L8������A�@pJ'䯖�F}�e�3ƀ�v���y��/I���{_�M�To���:���hZP��B�U�}�rVv�-� ౌJH�Y�(8�I��l�K���ֶ����������.����.^rt�w�U�p�S�r��=����9���I�L9��L�����l��I���cp;;.F�x��j�-D����K���kBTw�3n��}�������fkp_��B���7�w&��p?x^�k�w�.�V���>@ƨ �9@�	 S4���@z��d���-ۗD�i;��fU֠A��f�����"pN�ݙ}AA�����	�(15m�`WM�����4g6 �w�
|�
|�i�߃w����iD�9�@2�9��L?m���S&����*���Ă��Q:'�/6�]����+�U�vUh��\[�M�̞�{Xh�d�n>l��'�fC>a�ܠs�4VJ�S�㒶���L�fȧ�\<���6�蜣���0_�T�k�hZ��"|ҫ	6G��m�߄����3ys3=#��Ė7�)ǦXm��-����;��jn,�g╌c�P�W~�⻹�?�v�0��Wet*��ү3p��'9&�d�m��c�YN�\W�3{����.g������We����$<�1.�{`�/��ԃd�J�
�J�+���K(p�(�@3�B#���8�]g �!Ѭ�����-f6R�>��:��j�	f�	U3*c��G�����>�_�xl�s�b�߃(]ϖ��蛏���oJ�^(��|����n�/��b�g?����k�?(*���lar�Z/���ӏ
�Q��x����2v�#��z�ؐ/����Y��/_@��k��gw��xc`�Lf}�)�Y�.�Y�stF~l�`R�9E��kq}Bt���F�Ż��ǡ���=�^�GQ_�c�i�������ߖ���|�|��!���J�������y)9&ܽ��¤���Y�L�[���.���f��b$�'��a^DbA+��gPf�ew"��C�?��Y����-���G��T��!�����ޏ���Lit6ǣ|i�o}��J��և�-.�{,�K��$��p��M]n�x��^��"�?J9�í��C��������]&��T����x����r���
����O�@�=��`�#�L�2t�~���O�I[(C��!��w�As�P��K!���������/�0������ͭ%�v��"��٤�I#m�����Ჩ"�����QE�œaR�c�W�B��~s���U��FT�m+��
���)+М�Fg�T�iH-0C�;!��Ȝ��]��dE�K�9�D#��3G��Qz��)��$����&Gb����h#Qi#H��S�2Rd��ȡ8=ed���:�H?�"���|�:��O]$�"�D؅�u�d��g a|���"��x\�y�p����d�rI#4�y~���Q�(�H*��@^�A0�͐���"V�1+�ÉU��Ċ=}+��D���;�Z���a�ID~����{"�h���8�"�h�D��É��LK扟�?O�/��-��`$��žE�9��}ʸM�?��4��%��Ϸ\.gb��Ι8|��IE#g�բp&D��)���Y�c�%2��Ϫ�a�o �˕X" �ΐ ��Б$��#G���j�������r&&�)�����+_B!?�������IQ�����Y��J} �æ�ɑy� �}�"��B�0����D|���?�o�A#�a��1d���H�1J���O�U.C�M>�Go���Iߜӧ\	��29����8�}���p���pk4t��f�_�: ���H��1���o����3
�����y |��(|�g�k�R���X0LC�i@���n=��W�a;���pj��jPX�NE��u� ��d \�a�"sf�`���cDǖO�<���� ��������;�C�/k� y�R�	�l
Ͼ��eeBZ5:�隀Ov$+�LAB~�c=9��Q��g{%G��վ��v�lbH�FL�U�*<S��% �%��}�4�ђ��1�M!|��c,��,JEq$JE��Ra���Ow��)�^�=�s&��#J�d�G���a�_��?n�P�4~?��@B���wmy��G�s8��Ἠo�D�ȖP�ӄ�s�f�@�N ���@q�)
�b�^N��<���(B�=��|y����1��tK[��
��@��OO2�PR��"����Qy�[�Ru�Ċd�A��"#�S˄-B���Ҟ��*ͤm�P7-A����Et�����\H�M!(�|h�+�!jڡ���1��̷�3�{e�9Τ-ʣ����sKF-:�W����MnҴ�N��y��{���s��/l�	[�G���z�z���P�!�hژt��I_S�E�5�9��$��J����&X�.����  �G�o��� �gܡ��~Iq�͟Ǖ�q��ڴ�>��+��T���N$e�h��f}�X5�����sa��ֹ+�R�j�6�|��+� �Z�G�t)�� �z�%@eX�9M���g�� X���s���� M/�� \��9�X�5��J�{��r)����_��=���w�@&;����ϰK�G�m0�&<*zz����_b���Ҙ@�,B�O>D�F�B��q
�eR�(|#�z ��D3���FJ�����"�>���)��3b�y#�v;���Q�j��@K?��!�2a�\#RxIKጒVm��i]�k�EJ�����"K�%9����"�oIk��$\	�!�'��ִ��h1]ӂ{�����Z#���zrjJ� [jl]�q\�Iz����-�d�E��������T;�I5[XۅvJɣH䮖5�]5�-5I�a �V�w���~	b4�'��7����1�~�l�!î/P����>@�z�0.8��M������]v1�l8w]�~L;D��?�ƪ:���:Ɍ)��\�2sbO�2_,�R�/E�r�+�U���܍ݍՒ]��e�.�]�F�ٱOX�p����#���x/��b�u���qo.��Mn^'�I�������^8���nf���cr��Ȑ{BE�1���J�0#vhcw�(�������0F��]�������|�NW�rz_!ߴ���$������_h>�Y�NɠAIC�̭-��f��%V!i��S6F`yWx�!ـ�EFL�c�W�$d�}�V�&�Z̄+Q����vx�$)Y�C�?�O
I�����V�0
�>�B�(���K.��q�~�����-�ͧk>�ixY�ix��t��r�i8�^�.r���ȴ-���@4gM�����L�@ԸjX *��	�E��#���	/��}[�"�P��� �9e��2�uy��#�|����s%�6��QrjZOg�|��ߢ��P>h��E0" �d�w2�L������k١��(�F�;P���܁98"�Jn|��Zw�9v���u5t��!l�)=[B��Lp��S�C��%���6�p\� �Łs�*;|��|#4��$��By�v������.ཁP�,��eWb�om�ww,���_����ɞ	��P_�I'�3V���u�l�F?�:nO�Z�v��E��8>���,�<�]jh�Gh����~�+�ԽRM��%y̪�J��is��2t)%2K�(�^Yk�#����j��Wk/5��[a�a'�- 7��0..+���B�,SA�%�I��D���!h`'Xp�E�w���^�� ��%��X9�J�ϴ7S����a��M����@�x?_g-u���'ق"	�[x�sˁ�*�ϒl���K��Pu�F^��Xx@D���b���D���@�y/R��/A3����l�V�9nSC_>E���,��x^������M����ǃCUZ�����g�n7۫V@�'@W��
S��F[������z�uq���~���Hl�� ����Uܩ���틌���~�e�;�~�Kx���:�)4�Wi�^�_9�[J�ƞ��LBr~��a��'�$[�/9ؒ/�h���B3zt4�p�cv7L�+�cy/��C�����sN�@ck�U.
�"�Uh<����Q'4u���e"�6{X�d��
���&$~�Wo���Y@<���3�Ĳ!�l��q'��?-t�+�C����y�u��7����[g���F�hnN�>�)�xǺ"����$��A�@��S%�����P65!u*�H�{ZyK�n�_`C�9Pcq�/��hiG,���.��b���T�m���Ñ} �c�g_sE9���O���v-.Y�m=	5����s��M:�����[�G�,��{iO,oq�{Y4�7�
oF���w�y|������Zكk�x�aj�����|���mF�eX��}�(M�Jz?�z4��z�"�p��>d���������f� ����$�͡ѯ;��<6�/��A[O������`�n)8T
�mTV��>Y-�y�w��8I��������i���|�X��^Ѩ����jW����2���x>�y� 3�� N��S(7 �C���ç���z[tۯ0*�<?�R���\_�?��Cv��r2�؈��IQ��.�'��.�^j�����S8'�>.P� py��:�<U�z]�/��ߧp�T��Tv7�"ju�\�*�P�#�3��x���W� ����u�����#a=��>;\ �R���T(��\:�S���/�:a�a+�@a���v{��HH+�\���d�@��P��s�@���Ӟ´�9K#4=����"��)�K���L��ġ���y>|F;���yG����ɬpY���)BSqvM+p<�9&���<�S�1�3�qֻ���ψ'YW�$%�S0���������Ba��"�xA�����$�PE,2~U��c@� �"Wd#%P|NqM�Ɲ�DU��)�Ws�~|��x�'�� ���?�l!�\���	��ܠ�yދ�w��3r�<��Ta�=�Oe&��)�|�ӈ;qN>	��?�N);�oB�l�f{��䲍�=4�S�k��:P����I6x�X���d���l�	6�Z�)�(��|�R}Dq�-����M�? �*�(�Iy�D�Jq�·�z���}Aܙ�&�usm��<�|UR"��*�H� �1�\�t���2d�qsI�V|#��C��BV�Xx6�v����a}�y^�>�_8a��KA�����b� Y�dC����7����:�_��DJ��K���%ξ����~�[X�_v4_���J�<pP���A]��j���y�@�.r���6�}�=�I��� �7~��ٹ4N��@�-�~ l{�;���EԤ����}�Ӆ����X���S����~i/�_ٕ���h�&��Ɵ�@#z"�'y��ev�t (��2����,�ɸ)$96�I8���؛`�ݟ�M��rx>L&�R�^���B�gQ9�5݉B�E�r���I�3�6�W��f!�_���͌��d���`���hhAu�u.���rFOt;�$�/��R�kiʾ޷�����y����`�`z�V6w�D����	�c��W?xx:r�>`��?�*N(ʵ�
 <ߙ�#�׊��ޘ�րk��|��#�E���C&̨dM���:���Ʌ�6Ё�e:���)��������Q���-�[�-�������L�?�7�'��E�|a��G��{���f�u�>ӝ���y����1��� �I�jn�D�W�!�q�5�5^��|yS�o��~��Lҹl]��h�t��?!{�W����E�����������^�\���������/�׼�Z7;Ml���G��-bz�4�7G��^I�qv�{b���m@��c��6|��4�.�G�֮<J��P�
�&��]�#���}^Q3n�xGȓ�����S�m��b�=�B5��lǽn۹Ւ+��S�Q�Y���PE�M����J¬}l��ʬ�yۍ�~�f{ �˖��y6��P,��W���X
�ik�o(lv֙F_fI�m�����9\rx0�`�:�?%) ��.v�)lJ��h^i�+E �Lp�֯�&�����ox{�E�i-���ـ�Ÿ;C�-���ς-��d��~�@�XS��)�w;�Kp���qG����,���!�Yc-/v�ڼc��� Pc8.���>l��ة�}���aK�B�˯�^�Q�g7�d7:��X����EO����4t��&�i��WU7�	�Q�'.��M&�GG�
�6����6�w��2`=��y�K;X+qD%���U�`ؿ9E���ae�` _����u%am���\,�#�v(�є�}�x�����χ8+	�O�����_�c���?��������H��+7�@��I��Ct�����H�|�X}Fa��<�?����θ��P<*n)��u+�q�`x��T�p��+�~����u���)�8[�;��Ia� ��J����1���\3�8���z)	�Σxet��9���s�[�_O�0�����TJ﫼ʁ�	ˈT��!��r���AVj����$h[a��@�Wb�a���Ad�%)(�o-���
�l��P��٧�tޙ�H`o���Ɉ$B��sH���'�ol���a���0p?lr�֖^~��Bvխ�h�i��.Q|�ťlN���������'Ɲ����_À��t���aI���?�+����p�"�=��}J>jDd���J(E\���5{Z�whsa��Zb-��D_vi�h������*䴥�^�lZI��t�z��U���
�$�+w8��wë)e�9bw��Ÿ�PVs�P��@� ;����9.vV�\l�D"�V�92�a���u-o�6x[�Q[�`>���N$h����b�V�E��Z�98�{����9�ckE?@�kJ�d�����&W�#v�O��I�l��v����}�����<Yi;��i�L��́g��k���fִ�h"�@�����w�t�����*E��NȆ,>��ɆPnG6�.)�v:]���\�l�Q�ݣ\�D"�N��ƀ���l�(�fPF%�W��fk̑ٶ*>���&Wt�ٱ�i��wPŽ��r���v5��c�^�=R���e�$4��=-/,~R����P����yᰄ"Z|6���Ƌ[��QX�3�G�T�ˮ֣��q���C���C���%Z��hfm0��vtJ�9J�H�=YT�
���=iS5���$q���{Y��Mb��� �U���NO�΅t��G(�Geb5��SI;=�^a����]��aXԖ�/���\l$_�e=8O��=@�i��cw�i��`�p߁ңblN�P��WS���lJ�yW?w7c��zN��l��]=��TG9��kՏUQT�AQ�<8WW����0?��=8�;�iѠ'\�+��M�����e*Q&�H��-�
:�a�̕�3�U�,F���|�ÉRf���=]-Q�4�����4̠'�#�a���E�B��V;�\1^��q�O�]���Z�C`�]l���,.�����#򓋵8@zmGVM#1O�;	���Q�/*>ݑ���p�ZV�����?��Q���0P���W���qY:�R-ID�zZw�܎!+K����^eR(�$���u�G)���&e������	\��ˑ�Y�ռ4�y"=�;p�z^Z��M����R��X��{���+?�j����j��sW.E*��2��x!ݍ�AEΖ��C�BYۥ�,�Ԋ���ћ��fѢ���Cj����
�n�8�T�p(lW�1Bc&�Qs
���"ܶ n�s)���h\u+L��Dnk�z��s]-=,��33RKN���2Z�c��[�N�O�ʗR0��|���5��U �d\U�94����e>��"�N3�f��1S�� U���E�!e�p��w_���9y��~[|� ���uP|�m��[����X��}6��mO(�xAU��')0�?��)����4wEo�	D��*��x&�b�ė�ϒBE�Um�3Cs3II���;p�9��x` �i
?j����^	��Ʒ󵽕AoUߪ7�i��D��ߡ;srw��2���<�W�R�F�d�'	�О��(dX��$�k��tk�j�ڊ�<)�@?�#��d|I���i*G�����Fv6W7���4/��
w�S�B s$:$��E(W
�A@����V@:��?���V7z"�0Q������*�����I{�I��;2��Y���N��w?�GJc<�_�
�:�i;_*�Є�;
(A�R�n�w���q��W�F�Z�?6��:m?�96~g藈��<�1Ta�W�c֏���XN�,��)C0׍����z��Ll70;��2�k%��_��x��/p$�m$����j۶$�Ex[z�E�A�0�Cu�=%�h���R1�����~�<�8B���p�M�KP/?E�gؒ��s`��7:�oC�-���-q�s:ӕ]�:q1������I�+�aG�yjݬʄ�m7kG~��:Y��Pܮ�@�`�\a!�.G
���@_�J��Z)���H�e��J�7lHy>ɗZ�g%]�����J�򱱏��Q�q�d.���\�2I�����,t���7Hu�׵I_��0H�w�DⶔI��8h�v="c��:>,~
��<�z����;VaE�c��w:A��CO�[�B��~�V�~o�z	����(Agq������Dl�T�iTi-a,�Nh�Luu ���W�v{��:��><U��ƒ�����T�?ѮE�T)��vL�)B��oO*��(E�}��!=��t�hU��P�׹��3踒5�Q ����e'�����k��cي#P�c�\�P*K�S/:K?e�7�`��B�X�5��ޅA	&�� \���0����+w߳��qp�� w�m/):.����S�����Q���p0{e�u'��>1傌�I�W�Τ���0�b�l��"S.��X��a��j�gs��0�t����5��M�Y;�`{T�^~%���.>������R�)\p��>� �ck pO��������9��rV#2Q�Gq���o��Q)~lD?���'�lV�0̓d"Qj���G�Nۇ� �l_�����:��-��o��d5�p���z�!�ވq�]�b�������[�-7Ae����-��}6���>�I5��nh���'��^a�'4��G�{�5�иW),lz�t��&A� �y���]Et����=�|��g��ȍ�A�������M�JP{�<�Ҙu���gӊ���1��~R`���e4��"x�q@���I�]dT���g����Ƴ��0�,1;:֙�)���	P>��"�e	�r�����,�Zy�'�u���H70V��-R�^�u�UIxqo߭���9<��N�+!0�_�[���5�U��1��1�m\�{ŗ��Wz����/��u*X��#����|���q۷���f(4�W�{���V�rm�{/���/��Ib���c�����:o���Y]z0.d�.a�����\�/��/��9�p˸��rg��p��Ĩ���١L<a���aqmF�j{i, ��e���_�|�z�{:rBS��{�+>Oz����˩�<�8b��Ҩ���D�&7������a)b���:��"0 �CK�]tU��	�D�H�fh%؃DcB;;iL�
�%#D�����얰:	i�����?����(
bB$	 PTdt�9"k�YA���{߫�������s���y���{���~W�Q̢Mt)qE��#\;a}-d��y4�S�Ә�����'���)")^͎�Mg��{�o�n�y�[��0�\����c ����W�h"� ���8L���n���t!���tQ�.�,�
���~*{�߽�W��́�s�'7��O�:c�GI��Ή�~�[˵v��[�\����Z�(�5O�Yx�u+���߇�=���+���7���>�����1��Q��3��ՙhI�v48��?�o�K8�&4�ψ��Ad'��G���~�(K��}���=�=Y���j�$HO�:7׆6��a���^ �7��צ��mS�������`9��
�%-�E)=�6]���{��E-_m&��D��֌_�v���������������b��_�_�M�vi��wv%���[�b�3~��f"~�x+~�������{g�7��lD����X�"���uJ��
���d�������D���$%���@�����Vyc���rq�#�O��~K�Wk�Kld�ġH���@�'%�Rl?��ZY��mȤ5�sD�E��yB����8HF�p/|��6�q ���n �S��V��D��W4��ą�Zs���~=��wЯ�+qpod]��.>�R�o���N�����B@����J�Aݛݡ�+Q�t����c*X��@x��t|�LU%�g��A4�<�h��k�g:|�L��C��7*��-�!'D��ߌB�f �.Ev��6��25�����'P�O!�AGg$tl���t�v�kpqi�W䏅n�^���Q����N� "�!Ŀ��$;N�uХf��]"O+��4:�D�Y僁h)�)�\JA��R���u(��vT]F�リ�T&�p���*���W=򃦉�J�U�Z�c\��-8�B�)/׾A��/�����tȖ�����&�޾��ݔ�QKl��K'��v��W[���F�WN[�X8�:$�)�.���? �W�簄���h�[\DQ]97 -�gxXA�S������RiS=�Ht���7",������^*1�U��A�d�_ Q�M'q�
��&{��[������@;�&�*]����!Y�|ӆs�:��=4�� ��ć���+@�f/T:f���ƙ�NѵėU�ȱ�z\���Qs�ɌG�4�I��T߆����Ys�I�n�Q�	���|��6�G��Y~��gy ��ھ�ݧ�Q ޅM��u,s��'C��b��ܒW"C?�eƠ9��-˂q"�M�\�V�@=�,��ۧ�|�������f1���%�&�N�E�8,�)иe+hQ0�&�zM��ѯ2��A�2d���߂p� �rޡ|%��1sFc�����������o�ux��8<j�f���D����%�@~���{��-Püu��*����i�Κ�ዶ�H�~1���eL'�!�7��c��S�M�E��[۹�#:�/aq,&)���p@U&
[��`��E*= ��#�6a�Z } �zۂzdx6,r'K���g�%}~�;�Ч�I�^R�K�]d>RV�q8�]_4��V��j5w�-4؋zц���\B��D�>!�o��z�_p�?3��!X���>��D뺷�q_�A֟�u���| *�(g�CҨ(�8i�\l�r��r۞��ci"Z��8`�y�Y�&�;��o�&�G�9�nO,D�����e�����H��Z![$�+�_���N�hf *Ź�Q��p
�"6�A8׮fB�`[��X�4y�0��e�����lⱋ�Ц�5S,H!o.��M:p�h-��d,Qeƛ${�xJv�lf�._���/��Φ��k���}�I\��}װB�[dh^	�ܾW]3��.�
��.���g7���	�Z����|&$oo6���ַ
���\|����̶�|�~O������ri�ǣ�ܷUcI�#�ϝ4x�eb�E�����o�G�¶Iv.<�+?�VY|4`~�"�h�����*�9���q"���������,w����_%6|�1A�饎���^���Ůx4f=O��X1��k�{ԣ�[�)��`i�{I=��Vt?�$�`͑GGN�{$_�����I��(Ρ��(�'D��?f�"j����H�R>���G<\�g홉�~���Ў�p���p��y�6�G�⫀��W?$q!\����Bp+(�hL�A��`��D�s�oӸ�K`�W�\/��"zn�h��:c���#��!�r�6�~������2���3����} �G����!��7��H8����0� ��.�"{`f7xEk�}�>���K�C�{;GQ)s�1�ٳM�B�4���C�s?L�P�(Cۏ9�x Y�8��F��A>����?מּ�Q�,�A��4�����z��(��]�`f������ǵ�w*-��A���Z�܂��%\fa�YN�)r�އM���s��?�-�!���f,���\�XNi�����W���f��ȍ��XM��L�*�m�Y�G<jU^�R�	-y����_v�-��wV���?�����a�~��c+��I��x��N����?֤�t�(����l7��5�%�&�3Aa�c<��.����(�NXQ>����� o��Î�2�S8̷�͐�mΥL���u.}��9%�gw�ݒb�x�J]v<�{%r��xj�g�qX�����	����5_��*r\l�a��R�2�W݈�xȆ�C6�4aU��~_�t�þX��nO7����5z�G��xx��������[��eH��F�a}��	�\M���	Nw���@!�a�=�"�k�T.����鉻�4�f�&(%�l���C9�?)��=ߩi��-m����_��^��{��)�����L�-	�h�;��V��OOw�<:��H�Ｑ��$7(��}���h琮��q�i�? 	���wF
5�'O`gx��\�-�ܹ1�yzs"عd[�7�ſ)7*�Z�.tE�Dz儿y���x�rn����i�[�k��)L��������-�>ű����>��mn�{�&����������ck�77n���O��$䒱5��5��{��M�ƴ24����6��-�kz.��7x>�b�� �aPn+��E�
ZrQ��z]�&�������H��`�+3�7��ނ�Ey�/-�ʉq�d$vT�{��nU^"Os�{��`�v1�ß7����[('��cCn�	�6I�= �3#4�9�� �c�>sL��|]�v�=dR��&��=����,��}n�r�,?�Oڒ�,���d����"�h9�rNH?��_�*�
J�M��J�~F��,am���H���J��ҏM�����gR����2�t�~M��������m̱I^:�Ů���Ƙ��H��jLW��i/��l�҅-��S����Q&_�i�I��wi�[#�����+��y#�,qi�Q����W��-!���a\зc(!%���}v�ir<��ؼhD���y��qZc2~8���X���nL"2�aY�1�c��:�!�t*g�YO�h���]s?^C��SI8�`_{��B*�
���~X�5���q�s�뿟��o7V[���j��m���� �\PL���V{�W���xy���¤o�����"������_ޅ!���Tߺ�`��/��Uې�o���G�[��ϛ��M�'n��_H�q~�>q��\��MaC���¬o����[�Y�f�PL�\Ԭd��^V2��\�G"&@J��-�l���<)������ؙp����b�P�(\1����İ��DGq�N�x'�,V��a��M�
��C���Et,W�r�|'�r��ήģGJt�j��,���r]?�ͤf����r�ZW�5��1>&�c��(�#|f�@xz�W$<��!fiWO�'��+�,�`Ee�l��<��N���t���㉲��W��Bv�v~�Sv�t��g�!��Ť�[Mڅ<��ZF^�x�]8��e��Xs��Ž�ْ�xU�d�~���5�oA���W�)܎ѴL�WhesL�߃\�;�/�~i��G��l���$Քg�nLh@Zj2 E~��q�I��h�m��[`ejE>�Ʌܕ������Q5[�Q6���*R51V�g���U�ܢ�K����S�޹g_��IP�lelH���\q���%u<l!�T�W�u�a�����G+e�s��8�>%P$K�VmyG�ֺR�2!tWYU>�Me��P	wT��j��2:'޺7ߐ����8�&G�\�ʵIn�l�|�������Fw1���VF���2�X�-�oPh������B��.��c}<�mQ�qўk��3�G�����
]��@g	&��M�^�u@�ou9L���ء�>�,�PSn�����Z�����U����vx�����IN���ǅO��duv#d}��7���_��(��F��^A_`������+?��H)��X	������ځ���6�z��a�gW�1H��}̽mV�F�\��b�w���%�����K�����4����l�m+-8^R4�Q�)E�� ��i7����������YE#���n���3�e�\�;Y1�RտwB�����/R��?i���s&�.d�,��R��P�a[}�L���ʈ����%,!��_4��\�@��p�U����E�J��sm�#�Yk�"���_��(UwB>+X>?�
=k>��|��|
�-������ឲ�m�8�&�8uw`3�(VϺخ�����)�|����I���Or���]���4R�M�S��q���d�׏�e��a�S�����r�O��q�"�� goJ��q9�4��`A+8R4�Q�<^e	�e�s� ��ۜ��Bt��|V��y���=`=��Y�a ?�m�4����0/��k�o��݁앻�D����gI�jenRn*�<S,������5��#)�.|l��﫭���Օ��I9�K��KQ�-HH�D�]�V��4���xP5�j�?s)�s���)�~�ij�o�^�?=�/I.a[�4Y��H����-3�b��Chx�����!vp1�F�8�JRx��#�*1EK O+�q�Z�3��X�A{���+��`��ǒW���49:L�+�u�g64He�a�k���H>��c�p�!����"��5��o�I	F��~A�M�;���߿fߣ�5��:k���fm�m���c��3D홯�cᢨ��M����
���2��i��G��n�PG��M��:�za�$7I�&1Ro�S�Gh/3�sXq}��YNI�lb%��w��\2.ć�_�<e�W^n�W>� ���9�Ӝ�NK�?t%��'-|�&�.H���zG���0mA2��b6vF��Y� ,ڝ��Ü�
��;4z�2PF��_B���R&4ث�O�/8^4P��d�j8#�@��_��� �V�H�&g��L$�ɼ��t�'ȥ�)� *�d.~�ێU���0���K��3j�;�F�M�2ɟcg{�Ŏᙨ@漆s�ի���w�m-Ћ_����Q�|͂��t��`S�Ҳm�i���HI�s�eD_)h���v;Y)�#���:J��P�P�=X��u4Y�t��D8"�MC��Il�,�[޶��r2c����ю�ޒ�~KPnV��Y6Q���g^�:ԛ�Q�V�G@cdf�]�Ƌ������R�j�{�7{�G� 3	�S�Mp�S�րAEO�E�]Sz&E�8_/���;E�(�2V��̘5sƴ���:9�����ѩx���x�4�u[�i�>73+��U-f�5��@��^��]��.wiU~�����_*}�29��W`k�`[W-O[�$�P^���]���[������,���PW���,O��my�h��Ǚ�g~4�}�W'��g���3II���ʥ����}�h%Q��I�ｮ����pL���b?�D�Pc�L�|��+�mQO���Y��h
�(wq��M�0O1�0����h�����	�C��W����(�ϋ�J�+3��a��=2�K�Zi�WE��ڥp����s��W̌��G���8��t,r�b��%=>�h�j��EnB����WoWe���aIT�5(+�(tQ��ApTTL4R|AGEE���Ѝ~���յڬܬ�6�_�i��.e/�km��Cd����e��s���;/~�������s��>�9�9�����&�zJ�����<�m<��gvf�]��o���>!���&�z����\Yw�Z�<��g�2�aNAG�]�h�=���Ų�n�r��6�_���6+I�����/	E�v�Ƹ=!T�H�K{���t�JQ��i�P���@��9<�]޷�4S�5�T�_J��:��r��]��O���4pg�_Ç��(��a�G��|�@�������+t�Ǜ��{����a��ֻ���[��-��/����������'���I���t�����z����u�?���_���������W%)��C����zN����E�xz��ߗ*��;K��n}���v���R���y�����J[�ϯ�[�믏����s�_�������>s���j�۟>'�����߫�W^�b#C��*hKU6.�+���gw*��p0h=��S(8����&���h���tY��"�)�x�-y��29�k�CQ��m&��S��٠���~�9ތ��}xU1
�Du�6���%l�#�P��PY8b&Gz��1�m��jrE��nSI�@�x��mmyr�2�Ą��:�</��aSnEV����/��;��%h$�|�����2�/u��֧�� �.�m��-<?��ƫ�Xօ�um�a�)�0+�1�����EA��}5�`ӣ�d8��_�<���'8�+�g��x��~#$~�~�z����A�/%t#36NІ����%�����W�>!l�JI���_UNzu�O�}(iC�L����!�Եda#/U��H�1�|=��n2�.e W��c��3e=�_A��g`e#B�S1ML���C��r��q׮�y��w�����8��̭�?R��X	�P��-��e`w2f�Z_(�%k���8�Uk]H��:TC	C��z&�/-��5��vo(GP���� KC��F�nD�>���ύ
n��G��A��8�!���Nq5��7x/K���(��|Ҷ��}�C���0"�rD.�{�GfNI���NiH�J^�%IK�%�q�����̖�f��kT7�?����)���x�B`��z8���\�V�ߓF�AڳKm8�h.�n�Lb��Lbw�Lb�J*%�3��[ 7�_�E��G Xޛo�k�f���6����	�>Zf=���+�qbB�&����	ّ%�o! ��m�x76G��Lp#د��<���p5/7����0Jfq�fL��\�����)�7���W���v�6�Պ�?�|U�O��B��+r}��p�����E����>�������R�eij���l�e:����}���J?x�������%7@?85K�D͖��g�_?�;_�<2K�<^(�6J�_��~ �ۧ�q��~�����gI���~��@[?��7Z?��g{��ܙz�����~�>����ڳ���/��g�����Ͽ���%������{�+��E����	�'�Ak��4��-0�"�[�+��w��?Z;'3�\�u��+)N�O��Bd��Z��q�/!:�+��3��*j�(���X"���o䦕a�hF��$DJ�Ec �8b��Ȧ�ôT[�hCQ�������/?O�t̺	���������J�O��^ ���R�W��GA�� ���{X�0�,$U�6�:��P䙇�B���vJ��Îۚ}��`�VI�p;o������Rc��l�G!�F}�S� HH-�Ǆ��X3Z�]��D�?�0�/���T�jt�]�l�nHf;I9<Hy;�)P��/i~�i滳k�H\�&�����-8�<+vq�S�hRF0�섣�e���&M�\G���f�*Ƈ��M�ĉ�]�
��A]�ji�[B�MvL��L�"���\�>�}_���3�������a�������?V+�k4(�)���α����p)��ϟ$��p)��{$��=����h����[5wz{�MIm������xC	��3P��p��#h���l.��W���=4������=t��|"\:�]#V���蟄�z���N3�aT�<��?���o�A3����tZ{CH�1�����.���9T ^���i�!�6��L!��sUt<���y�)h�ȃZͦ��'��嵱�@�}�5h��	���9����2Ci�a��ĵ~?џ�~J������E!���d��G��g�\��y ^�~423�X����7h�O�9K�g��7N���PFsZ������إd�	v&��š����&�@#7�i��e��e��k>Y�*��&�jވ�܀�q�hF �
��Z(
(S����|U���-�~w�J[}�unJ��JV�+,��S�� H��t��Б�C�	���_O�3��mZC�H=M��w)1Qk�t���ӡ!6�Xv��}Ds���9�{��,��1���,D�3�.��h�W	�<�Uo�*�Tɋ��c�8��'V�wMK�;�#M�$̶��ζ/&J�W�r-����t�d���r-G*���RIߜ+�t�\�q��Ƌ n�.*Fa��߬���]

�b��/h��Nr-��/`�To,`�TC��AWP*{8��?����6b�(5�@��!A�y1)�qT���e�iG��YZ�g$�n���D`�4���l3�TR���5���;=��N^E�P�<��?B���E���Vq�$+[��۳o��"g��F��L����?r$��o������3S�)X�
�&,��l�bZ�7/��L#2���V��{}>5�p � ˚#�7�@�����f�AG�@�8����ǜ��,��$���'�D��}�,��i���+��%�EeA���������0�}��(�?�8��#�3�\�iԎ.hw%���t)��w�Um�-鱍a���������.�����F�Y�?���IN�.KPΞ:�W�`P"ﰚ�jhe���B�S����짭����
��5*��$��TP�B��oArj,�-��*fɱm���(���]�����v{��F��[�t��FmR.�`�
$�Gv$nI�>�6Z��ZWN�)+�:�?R�O�nV��(�>�45V}9^b�
�H�U�9c�g9��*8�J��{K��̪��X��*@���Ŋ�J���E~�hp^�T�آn���4ԍ+���Jl�Ρ;$�q'm���i���0��8�~I1~�&ͅ �^�p��b�&�~(�#<#6����OX�P�xr���j�E�AZ��Q7�\�C�U�P����f�4S~bQ�P�!��:���M��B~����8lN����z9MP0T0'�7,9�u�F��)��Ȓ�<�ၓ%�@��V��M�5���B�q�:-�C���䯼���� ����V�4a�]2Zj����6�����S�4�K_f���n�e����B�<��{�B8�4u?�V�rS.��xQ��:Faw��"��7I��}ݗ�[�����?�J���J�i9V����]�m�P�2G�� _�.�#�2��+B	<�D5��bkB�җ��C Ιɰb�7LԐ�ldy&�߃H�E���`1C���� PYj�z�駼fߪD�.%ү
�"B��T"3��LD�Ϯ[�D]�F��/&21�鍤?�^��x"�#���Q�B�����]ֶ;U���G%*_7	O�h �)z�� ǉ���!#U�h�#�"�&r�(�E�ž	]T`�GkuQ�݅�vp�T�{H���k�ڃI5�J��sݰ	��ͅ?O`R=��I��"�T�N`��N�TϏRHu$emk�.k���b���R��Aȳs4 ���zB�M��JtصW�ch/��5z�c/���[�'�6�`�ۤ�}�A�fc�dC�rg��l]����',J]JU��5���C��Yp�A��8�`�E��zQ��\/���Q~a'̒'&4ʱ�8���Q�q�rܘϦ�m���P5`N��84(�s�沛�Wku>��+��3���x]^�ܫ�ϋ�C�
�����%��-��"$�T��E$��^��L�Ƌt;����l���
QD�w�k�Q�=�k�x R�"T��Zq��w�V�,��Ӵ�*L�Á§�[�b�eh�ۆ�I{����j�J6�V��t��R��h$G��8+�'��#���+�y�8]aM��;����bez���Y�f�;�KQfk����4�HƏ��R����b�9Af��D�7evh<ʬ$KCf�#��MH���m��4�]!۱2��:~�ाM_wg��D%�c�C���`��+$rW��ѥ+�7��$�"rxK��%�|?�����D��J�n��{ݤ��M"�!�P"��Ր��#�FB���[�Ii���$2s.[�&�U	g����ob�0�^�fd(���g�8VW)*a<Օq��k+k������h��R�x�T
�E�v�\՜|���j�c��W���&�+��:��5G���F�ۘ��fT/dR�����"ō1��0s&���L�#�Kq-�M�i� �k�C��05��[��Vqhq����U}T�}��(�!�[v��/�3"�yЩ�O%��B��$��͢�O&��$�۰Z�+��D��z�I�~_lw�i��G^$�组0u�?�6���E��6ta�����&r��?�+
h��,��q�+$=w�ѳ�C��!���Є����{�p�v5�+CV��q�kar	Oi(��͸:����(�����Gk���>T
�n��sѨ��:�.�?�y�4?��wC����-JQ��9 <=Zh�l���Ӣ��\h��b��k�>�U@�ܙq��3Z  �v:}�;4 =L��Cd��R^g4����
۵���hsg(�٭�=���*`��u�ϛt�ͽ����@�d�M*�<�p��bP��z��x��5�>�x�,��L�,��Xj��|��#a騏������ޯ~�������T���$ڿ:u�����#5�GuX���bg�;	�O�t���KH\'���e�
h���Us�/7r7y�I�e��$_53�ϛ��qh)`iѐ&�-�D� d�Gh@F���wK!+�6��O�e��+����.f�C����_������!JM�ϑ���a�����5p�@�Hq�W�mp��FD��_������Q��h$r�o�Z�)n��}��g�L!tOF0�24���`�K
�=bG�#0��-~R`Q�ΰ�4�aq�>�߄3���w����E�����>	��������;�X�*v����Q��g���t�_��OM��|��&Y'�\g���>aX��C-��� )}��bM:��3��F���<ӟ������[5���jc�q��C�_i8<�8l(���u6���&��_�`���i�����t�}BÄ�ڶ�?ܯ4���4Մud�;&��WC5ƻǻk�t��Ŏz�iO������b`ý6���T矱*�M:�|��X-R\e�Cr�����$��y��D���6�����F����t����Q�
���ƛ�� n\m��w��)�!��Fܿs{�lC�y]�� ��Hkf�yz���)�i��T3 �3�ƿ� ���r�L(X
Jա_����n!�M�:�`,7g�R#W��ȍ����F�*�++3r�䯁�=M�~���^i�bV9y���1rn�O�N���B���F�˃Fn�C�*#g^G�����F�6�6��7ri�\���\*��I�|�l�%�qL}���`�;�Y02S�Y|�odb(��E���P�ea���_E͕4����]��v�P���QLo��ȗ�8���O�F^@l�3�]�R�,�em4<˱�'�>=��+�r�3�2(?hJfC��I��'�>�YG�"Z$T����Z��T��FOp�E�U75��ь�� hu����מ@�N�#`�+ �YJ/ �CK�]{tTչ���3N�dĀ��+�<�!r	�
T�PZW\ƒXz�0	pz��W]��,zU�xi|y�G�Y�V
VO�#�s��}��9�����G&��>�����~?ԫ���n��YRs���#��xz?�Z������F�����o�˿ �	�.HI�P�Y��ge�gG�i0���_�1i�
�A<^v�a�k������<����IϽg~B=w��~р_�x%�z<�r�\:���Ug=��܌��'^}�Ic�����vߦ�t �ɝ^	rr'ĉ�)��� �ϕkp1)�$U��G7J��W������>R���S*'0��*����Ѵ="~�Y�_�j�k�80�k��Ysmw�?��㳪᎔���>P��}��D���'#�jdH���k�!b���N�t�s�+�s�}s�zK���&����ªH��F.k%�����2��:�����1l����Wx��w��>U$2�qѠS���=���˹-��t�:��Ĭ	,����T��.K�'�	;�G�λ�z�gv\�����J�GX|ӿM�p%�ɂz��x�_z�j����ڵ���~	�95%�?����O�ᢎ�}�K:(F���W������8��0x��)��C�ɵ*j���)}�y�ZXS_m�Sl���|�6>�U�3�#���,��+Tᦼ�ŧ8��Χ��ߋ7�|������XVl��������P��e���y��%�f�O������V�l�V�����\���þ���iX�ҷ�������,�ʾz~��3��uE��z�$^~���s��������{qqP{l1W�ޏ�P�/ _��*J0���'`q.���Ƈ��� �.)TY���h��[ش�Sml�����YA.N	ez��� N��>p�z��PA��N$R.����.�W��Z�
#?�\�ơ�=�T'�7" ��X��3aA	��\�����B�:�$�%������b:��]O���S�*�&����	W���{/\�����߸��������)>�Z��X;Q��a1�Au}x�1��,��040��GVZP�`z��q��P˒�(̑rRn���?� ڡ��`	��T��r�X���%�^��ïn���[]N^V�6��%��,�W�g=�h���WK�K���4筸l*Ϳ`iN���kS�+ ��^-��wocx!�s���%l�`�X,�����=i�>;	�y�9�5����T���x�.Z��K��x����O�g�P�����o�3�AI3����f䔲��m%Ĺ��3=l��Fd�$t2ŷ�O-llI^��Z�HOI%^U���T��S]ੴ�|��?\_��G���d���Y���ꦱ�C�r.lA�ڒ.�l�kp���,�Vm��b�M}�Id���	��U�>����}`-�`�i�~w�[��^O*AF��9�9���㉧�nB��_������iSv{`�
Hs�?M6�g��� �Ri�A8N����AR������]�tv=�Ji£�Wg=��(�zЁ1��}:Z`��:�>��7��о^���xO揲y A&�zs+�ĕ�")#���HcLk���w�?��Ӻc��:��I�.���U�I�/�}=
�z�a�s�\j�e�w�ꤞێ�/�R�kSm���<]#iM�o�s�H\�B6��4O�5�cN�o���H�g�
%�&�'��~��FU؛���+U���x�*4��bU؇G��*�7���X�jq1��Cs12���~��[	������!y�&�S�ۯN�0\��ٵJ�CU�s�o=�����.���-ވRW�����[k�Ж�V�1���yX��'o�(u��ʘ4-�3�V�{̛�A5/�ڵǔ/Wb4�fnQ�B�
��ROx5j
���?�M/l�A��,V�<�Ar�F���>�D�W���k�lPg��Ừs�$)Y��J�Se�S�5�G��ew�5)��Ϳ�uT\쐆C@`ō�^n0�&&��U�`����wW��W���P�+�G=[-�^o�1��[��7䥦�u3���E~l�N �c�:�pGV��&�d�&�\H剬�d@���7���"�k�;dM_HzJ�'��~2��%��-��H��>ؑ�埧��mr%J؆	��Xͭ��'����D/��0$IUN��лԟĹ�8�e?`���)�ǈr)�5��P{��v`������5�z�\�f�q��^�N�_��$���)�g84ٯPtj^UP�?'(���#��'r,}&{�7*o�Y����Vx�&����s֛��b��S�;A�ɬ���2�A}1�u��Mݻ<A?�S�q}����ž��锾Xh}<�''���e&�ᛀ�h�s�4�<��	�]z̪E��E�/�Q�ȓnG�X�^/�y���I��p��"n��K�I�tdԏi*#��%VUV �wNJz�ڑi���e�wcZ��C4� ���Y%C@�!�թ��"	��2���d�A	�t�����|b�����ev}���[8�E��fj�\�tO<�(L��_�8��.Op�_A~�Y4=�h���`���{�#��1q��|�����/V,6�b5*jT�A�@�nw�?Ө�
���2!)���?%�IYV�"V��a(d�|�M��_g�%�n$����	��R���E[�Xc!�mMr��~%����$W��$M!�n���E�=�+�m�#��K�kE�lG�*_��b��M�wtͩJ�"��󵤲_/�v��0Mo�{�t���Mu���j��K|��N�������Tw�#��A�$އ�� ���6c�%\�w��7(��a�lF6/�h���Meq>�Ykʁy�+:
J�7��C�J��}�#
y�������+I�U#a�OM�bn�	;ø��2SAo�[J��b��T*fʩO�� ��:��xY�'�`�`����P=z@���s�>��z���6=H�̺��C�D�뼆��ѯ��v�>�:���O�`|�L��/6����Y��N�ُX6ĸ�~*ݤ?�X����Q�\�MlcK������co�8�)���ɟ�����~��'~r��?=O�_�����>g���>��������i�R;#�,��D>s#�e�����jo��9��<";\}�FIQ��T��]����p�����p7�B��k_��7��a�b+�������G+�k왩�<��m݇w�=C��H�˵Lv�;�j��p����͆�L4���+M%��V�y���ib?�9��m�páJ��G�Ua��û�l�.�m?���c>��'�|j�O���'�]��l[�^�	�e���^U������Y{��Gwe\%{� ��̋1����'Tal�^�\���jF�A�R(.i 
2�I")=r� �u���cr����҇�����bn[2�n߂�D�|�fߢ��.�T�N�wҾէ@�o5�RmQ�xbd8�Ⱦ�1�	D��a+�m�aef���t4Q)�?��U�Gi��AX��r.�Uɴ�x��x������Ŧ0�)�A+�
��|9`��[��=f1��[�h��3������g��1.
�V�b=�֐T��
�)�l���U؋���l��M�*p��IB+ !X"u����W��#�:�1�'� �4�<D3��e���;؎�
���E�8~�X�z�'G��"��) �F8����7hS]�˱u��bVJ7�N�h6�f:U�wR6}�`���T���T/�z�?������S�K�iD7���ǳ��r�<<����ǳ-������j�9�ٰf�-��W�����OŲ�y�	@b���۬�÷��gW#mٳK�ߢ��Z�ˈ��ӊ�����T�����^��.�xG忂r��m��q �e"��e�1�I9�?��g�f�B��]��"ty�Йz઻�A�'�0]c�bŁH\
�%���n��2ُ�|�}ŦZ�oq�,e���*��xғ��E�c�أ�f�8t����\Ww���'Z�S^�I�Vܽ�"(cya�	�^z�����x�l����Jb�!�B��E��<��Lya>��J��M%ώ�����Q�u��dl��>�gߦ ��UpM�U����JJ��7�9w_V�51n,��@�Av��7�d��T� ��"���d��g�B䌀"��_l%LE��8��Ш�0!% ~W)ȱu��Fh�a�]��AAC8��q^��
ݺ�j$Ŭ�:�r>�tn��P��`y�V��yV~�����%����Y�W���l��FD��?7��My�����������a�sE�ȱ
m�-��]����X\AoH�t�?��NV����D߀Ui{�o�j,��?
��qk��� ��D`���zQ���0L��~���MO�em��k?�pẴ�l��d6�餉H���E�#�Q��p@�\ɄAy
�,g!^���k�ؑ�p��|pI����:�r�?�����Im��%�9Y_[@Nٟ9��p��30�dF�{��]k�><����N�Uk6Yլw�)��=Ҧ�Sr:<O�x[ {�-O6����6�e6f�ڲ�s;�a��7S4��ț1���|0�br�M�^�oy�d΢{����nby��~Ƶ���UD3r�GcP��3r.�qYJ�^襸KqC��v��:!By��u�M
���b�:�x��N�z�(OP'D�E�T'D�'�b�9�����6����[
m?��â|j~W\�T ��Z�l@�׳�H*~F]��_��j�{N��@���>��܃az!s��̉R���5;P�̙rΘ9^=s�0s��2�n8'��n��}L�_�C�d�|\Z��e�R�%�����b4urI����4��A��?�߁��G���1���6���Ym�L��"�ҴSc�ԤJ=Z��եC�KiI�斂q@�x(j?�X>{��-p�41�a�,��AIj�0ʮ��:����`>zD�t��"r��ç��.��<��,��6h�m�%D�(FֳVY��Z�N?y���p������W����ڴ��ܒ���=c�6>�ڈ	����7���U���,6��c�!>ͩ�8ȰQ+�⃜���g�9�zn�ށ�Jz�xzn\���о�cن��;��n�_{ǎ�v{�y��nĮ�[�F|P�;>�|n<����6�����󧅈�����Î\Z����dB$���Ic%�/��D{|�fje}����h:�_�#W�/�)J�Ed���ls����y,�<�Kd�q��<���e/�������(G�:K`ˉUU�i��+�&=�P8�����[ȼsE �tc
��8���]��_�H�I�b;G��_�m�J�z"O�d[�VA9�IW1ZV!J�^�oy[�������:��L*��m*���P�Zm��p�ªY���I������x�'�b ��07���ʌ����E��D��_P�g��-��>g�O�;������ki�������'�?�ap�,J�d�֣���@�ct������iW�����m3�g����:w��賛�w�=��J��<�W��Ў0��\nt-�av��fË���P��B���I�"�-����'��~��lǳ��p�' � �&_��@L��H��������ǷB\@����_�Q��[���,������ڞU�tG<��'��7aIv����ĒJ6bI�����x��T�� á���1+'(ω��h_��x������7�+j_#|��>������{�$�:����^���]{��tؿ+#	�d[���wMi�]�]O8���\v|���G;��Z��� f��
f�@���%�f����!��G3,%C��S�8�Ā8�!�E����q
;�N!ۊS�	0�x����q$J����cJ�9�'����k���5���+��������>�?/ �� �� � �p��PE될Ƒ��Bİŀ/��@�r�Ǆ1�#w;!���[� ��/;�r~�p��`�����^d�z��w�MTt�_��U�7���P�Qy	��Ó�x2�NH�b&����p=��ڰkx�W�F�B��pE�B�E.`9����:�
��/�|:JG��K-�����s������:�K��H�?�����W@ ����xX�
�0޴�Kb���8��x��ގ����G�O���sS�9�ۛ���n�no��"Hϲ�.��Ex�uĿq'��WjcY�U�J�B���{��T>�G�+V4"ͧ�>u�>/!:�>����B���XI�X���҆=�\Ɗ���(Ǧtc�ayQ\7�Ք��l�CT6l� �U�['�`�Wj��s� l�e��ʜ��tָ�r��х�^�)�A��a����]{tTչ?��1��Ճ�e`�i����xW'e������@�W��E��bX$K*�$^��ZP���*W�P�� )y$<��#�G %���Z5`������LfB��+���g����������~#�ӌ���kѱu�[�;�ѱ5����&����H�2�d6��tI�?$y�L%W�m�:P�SS���T�_U�V�-E�v�~�Hl�Q�g���i��T�9�(�a�'��f7Zy��%��/� %��!�<��Pqh/�+Y�����I^�awֵR�,F��g]�w4rO!��)��]0����j-��Y2m�j�l��6c�B�̸�&�>�k�>��&j�3�ڧ������=��W������Ѧmo��}~ަT��3����M�>��d��$�G�_�����s��t��3���;�螯�jx~�}~�Z��k�;O��Æ�!�����Io����dc�h�w8(.!_�,�|=&Df��y��NG����J}��y��*�U���t�a���=�qW6�c�D�l�0�d6�{�R�	F��#%�`5��6#��Ŗ|��¨���5n�Y�H6�~��~�C�8IP��->N^W�'��mY�@�l�N6��e?�E9u�_��p�BH�;11�\�p�j�G��kF��-��2�Ŕ�8���
���+v_�@C�~�YP�F��-�!ݯ�����a����Aq7|�KFRe�K�D�CΖ�P��θA������0���u�r�{w`��2�a	�w�K�O�b��ȕ)����0t;�����A�o�1��I� �����1s�'�T�& �&mrs�'G����z�cMI�/������]�p}J �Ǒ�����Ud��O!|����ƿ�j�_W��l�#�D]������Z��yq����k-0��A��Xz��>�pd>Ɖba�����2�A6� �٤-�N�
�nT��A�EL�T�����%s@[/�.�s��ᝃ��û+��}�����4�Z�5�P�=U�.�'��0�4Q���5n����
�]L�����j&3�q��J�z�jt����J�����5�ǿ��P���i'ۇ�S,�U�C�cw��;�� ��T4��nĖE�e[�7!QB>�Y�O�'ة̺�a֥�K	��8�ΰ�G�d���'����B�]0�be���͙aT�G��U��-�Q
A4n��-m�T97[�q��I�~ �`?#i)��0���O�����/uޡb����q�a;4L�'y�f�^|�l`>9�).*,�' B��0(A,$�� �#������2�������@���ܬ�p�!�p7����U�UD;�8��K (���c�v�wӓN��N��d�/͟1c�ޞU�{�gy���M̞�5ڳ|{��'{��ʞE��lI������s}�u�سFN1۳�_��It/S$�A�Z�nN���K>f�b�]-����I�_��7�č�ݕb���S�}~�iE>����4�8�7�SW(�T���e�I��5|������iѵ�s�uU�F�� �����C �U�߁��Hߩa�.@hm���H'X����!�8{��
Q�R׽�c,�/���2x&B�R�o�v������Zp�l� U(3N���GxK7�"���'�ְ��FO�39�5��q���=��ܞ��s��1߱�6�å������ՙP��GxNC�6Ғ6�,@i�xmZ@<��i؆��}GAޛ�Se0%ۑ��4�&�G4廔���E�E=p�f�C�h(M���ClaE7>}�"#����u�&N�����?ʛT��v�'X_,D�ol�v�='�nt�e�;]�ݹ��`�T�3e�CЃ��*�=�����}��T���Q\���ӯǯ}��c|�]�9%�%g�G�!eJs���u�]�!�h����f=����c~����"�����z_r��5�n|����b;g�D�g3!�n!{��D �,IZ�Pa:�A4u�5��M���]�Πv�m���l�e���FWJ��.�_������~֤[��M����x=�f�5B���V�L��ydQF��	َ8F�9ߡ�0��t��U��9Ƈ�UM�	����}on�yJ�?�������яp=�1���1��܃L>W�F��X�vh���/�=��P���m�2�[�v0�f����|�*��,0�U�#o5"}��,!:��y1��3�Iv��-6�����Olȭ���A���SH�|@�q5��ԭh������M�uC�3�ĕ�3Q]_�p	`���ӡEuD�E��<8Ԗey��@g�]�J�L�N����b�2�a>�I�8<��Ƞ��B��fJW�;�xt�Qh�k�e3d�F���_^c<�5 �1^� {KިxX��W���/�T�x,��4��cr��щ��pf{��G�~�3�fL������F���.�d$�x��%~��>t|���	�!W{��<�X||�������($�a�����8MX�����Q��b����6$�ŕ��},ŖLN�-I�h��~>���_ZaM��V�ǹL���8v�qQ,=���p�o� ��x�0;(�!�� 6�	\L�`�,�R��E��!�\��s�I=�t��8��a]�_�_�R��K3���^W��5�e�2������4�9lf`��ދ8�UD���6�&8M5�j�ޅ��4�D[͓X������ʠy�8T$��[3���qU�a�b��pj�8,}������r��4">������A������1I'g�8�Z=<úV&<�CF<�G�Q�I�5��Z�`ǳ�M�$�!DJ<q�� ��qB��*
?wUGmZ��� �y����m��ݵ�����/�Q=Q���b�"��I��p���U�k�opL\:"�)���P�AϵC���S�E�b��п	%�Z�!��D�@<_0
��(�_'�A�	ۗ�XZ�E{��.2���k ��辚㯐�
����x�M����*Q�@��կC^������_�)~�
2-a�&����Ӕ0�D*;C�
�{�9Q]�2\�z	ĩހ�4)�y��Ƌ�ES1T^S���MGV��d��*n�t�7�K�a�D̃�V'_U^ KB���l?ڶKo_ySw�~􊁿р?0>oexC�c^�p�!���`��_=�����u=�:�:��-���ڗ;Q^��=r� ��H ���0����}O������Ƶ@ʌ%%J���m�S�|m%�d~�6�)u�4rJ�d���y�N����g[&����X�$Hs�Gp��l��-�Kyd��?.h��ġ��W'�l��<����|�9��v���۾��������"��1�����t�M�#?K��R(\�3G�q����<��|A���|�aKJ�0�&-p�I �2ۃ�zU�{7t�h*�{�:Zw�(ux��qT+uT�,u����y��7�D�xDX�����b?,��1iN�d]��`V�1�1�����T�K`��K).Y�i�@���Rp�uy��y~ƟO�C�'3?�II�3:L���Z�3J�`�b�]�3;�R�e��팁�5��q><��i۔��caX*¸p�<���S�=�i����J���{8�%��xd����ƫn_��	2� ��M�5N�8��1~B|�F�|v��J�}��P����8�G�h�r')-�����>�^//2�#!kq��eM5���t��!����@���(C��F� ����9.Q%������׺q	�!�_u�:�ѣ&��2��?�("��Cr�CZ*���@Vw�Y��XG���1�H��+4�}��ﶗ�ed�Lv�����#o$9c��4�ί���BC��L/\R�͵<�Q�N��3Bx��"9�_��ɭ�����r�nZ~����_��F#)+;?{c|�v���K���M+ع���kn���T��ZH��{�*Qd�0��+$���,�]����?���M�G^q��:>�f��_Dq�# �%�B�a��Yi���c�E��dRf�x"7�0�GՕ�V�Y�*��$�����? �7���xp�-��%��'[z�������W��������D:^�����V^�I��j�o��u#Fo�����|��[���X�@Vm��w��NE>Ο��q�A>��>�g��J4�p%=�ÕX�Õ ?��ے�g.]�[{�&�Sm�5��t�m�g��/��H�g��_k�l�o�g6����7�	n��)����4���`�E�ʠDUdJ� ��Te�M�{#�}R���o=ގ�Tm��.��/ !K��f����t�x]ׇ�Z�f�A��?X���V{b�NP�����d�A��Z�$o��AsT��8�Z{M��ۨ6a��IA�w%L�����ʍZ-��9���.��'nk���;�eE�I��Bu�<�~g�S���5Q�0-?�h>Q1�p�#��4-�k*�1�G9������X'?P3Y&��t��y��w:�}��`��n�ˡ  `�d����F(R��4@�P��c��e�@�4��NFMF!K1'Ĺ��U��R�pxėva�/��&]�s�w%�}��,Q�l/��.�a�[|M%�Z�f������<�TI~rŬ�/�iz�	_9Y�x�F.,���*���Pcdl�cz��N���%#�.�T:�V��!z|L�6��U2+�_JI�Y� ����P�O�Y*�C��d��#�벴{Z����g�f���GȫL��{�W>j���mIJ�ٛx�Z�݋)!k)��.��6�ˑv��45T�O8�ʵ�W���Tr�޿1~��1�bc�dq����O�m,0��q���3
��@3^21��l>�d�# R���#��pUG��F��ܛ���E1�c�"d&��P�$5h�"���*v�?�6�P����@���2Hv7*I���a��~K~U��]�j�`갹��\Z�qa��']�*l�rn,�13a�Ԛ�޲3��A���KK��VE�VK�+4_My���ט��tvf\*��^̀�jJ��V�Hd�s��[0~?O���d�ʄ<���k����S�^�lY��%���n����^�n�+�I�R2�Y̵l�����	�GJe����{�4�k���ߎ�1W�\ܐDk��8�"�0�"�=R�L'�7�tK"�,�������U��ʹ�U��B� _;�!�9d���3C_�@��/9Pc^� �]����!�H��S��ߕ�J��*N����I�,È�����ׅ>���@���Ð�?�^+b�("f�a���ih���W�������8D��}�,��b���/���C�_��E�����C���)�xS��/<�Ǖ� �e�d�M�d���d�ѩ���:���\A��h��XO���<�,��G�"����!�{nƑ�k�Fy�����APC�����l���Y��G=N��j�Lk}{bE����@K\i8����2���b�J�Y�����bF�ե���	�.gm� �v͝C�].U�%=[�����J�ĳ��󁴼�<��Z����$�v$��a�/ �CK�]{|Ŗ��N�ݨ q�j.ΐ	t@x\��J��BVX3�3<�$&cg$�+�hT��g��eA��}A�������l�S�=����庿�?�����8]u�s�s}�@�Ӫ,}/�� ��V&�==��߆?�d���)H|�/n����E n6�k�g����%��񁤶�{Oaʓ���Q?������_|xA���u�E/r�x�������}ϧ*����}�T�7g�ףτ��M{�kj�@D��v�bR��;�A\~n�9�D�H0��w��a!�m'Ɯm��覔&��){:��Ι8~G�:~�A�^۠�!�*~zm�ryC�a�����~H���=���D3�<����~��?4�����d&���]��\r���o@*��s�+$[��Rx���S�o&���;?@�p���%��*+��f�&]��Ố�I>�Ӑ�?(���Y�X��e�<O���)@�Q�H��<%W�O#��#�1�3�h��;��#�7;	b�;�2>R���Z���C%=k���k�f s�p#B�W�`��(��O��1v��U	�^�6]-b��;��A�,�_����U|���S|����`p�mt�͕ƻ�|�G���0[g��㝲Yw���j���,���Io�'5����~���P��m�l�7�7�s��>�ơ�s:����5�;UiP?S�"M��[�鵔��/��ǄC&���H��ۥWu�wj��Կ�:'�G��M����cՙ������}d������ܿ�6z��F!��=	|`;:1i����ԣ��Y�*�9oz��O�T�M��$P9�]�Q)M���qh��c(ɳV���S@~�ʶ�ImK�s[}Wg�O��Rs��t�A�Vy~?
&]@�N��7:L-t�<���D`�Ѽ&�������;h˸�L�����d���H�����\جUU4fmz��ט^��'ك�x�On��?�� �j��j1����chR�lb#�>���\��� &��k����q8�%�����>������	�U3�z0��ڣ�3�����> ��;���!�U�Ys)GV���xK���p#���f]	�?��@FP�vZq ;�z��0--&�\�j.C�a��i-pw���N��P[*F��D+��X�z��oc��0kN��xD�̥`#2�B����_s����4g��uv$"_P�ϼ����3�=�P<N^_W�����⵻8���Ҕ�;`���B�B�#��O�,(t2 l�I"T0# 3n�u�����07D�I9�Q0���^6�@Y�l8�92�q�ðˠ���0Ј��a��8�F��G��kQ������vO���;��I~'n��'���>���n��q(���[ �n��c���q`���I��>���؍p;�H����&�3�>�H����͢[Ȥ� ��"�����yI���@sw��jv�����oB���Dx]���k9������a�����j�_9�X�L86�&;���F2+�=q���,ݪ�b+�