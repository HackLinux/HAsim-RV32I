 
)UMvt�;%J?JCdx��x����P )
Gdt��h}���}���}��}+b�G;,C:)AsIR��R##IAA:Lr~��n\j���ڏ�f�y:3K��������յW9[������[266@@!\j��v9.GPRU4^x�7))Gdkt�v��\2?0)  4<)!j\j\&,%%9PWEk����tC0 8F$%	
	A��AK���m4F[Z8X[w�b$%;WnvbB82??--4'Urg�ԶxRgx<'34dCWbHWv�v2.w���ƿ8-Si 
34:�pp��oA:/RI3<x��JH���՜����t[F/)Gr�������ڵ�}$00t�����j9Q6@@@@jj�j&	;?;43<xx'7G4)?Pf�n���h.$8,88 8tW%,%2���}&+9,$2BW9$02d�d2%, 		
	p�uAK���FC���P)CCk��8	0Bjh2.$??%;UeR3����IK':Ig<C<HWvbb�\t$9w���h	��dF)<Ku��u�^AKRgK<o�i8,}���پ�}�h\S?4L�ÿ��ھ徏jjj	&9[�j����Q\jjjjj}j@.7C4))LUR<ZI:/<PX��n���9" PW�b-202\�է\.&$ $2228dG"% %		


g�3Ka��݇7C���X(<4d��B.MM\�j\&$%7NxU<R�ݳ�RIA//g<)NZv���Ͽd8vv�JW̚F:upuaAAR��A���8%H��վ����n@+\.	8��Ƶ���՜@j\j&&2bh���Ͱ���jj���j@!.0 0)<< 7<^I<Ui���k��2
Wt��9!99MMn����6!&!!!%2%%B8$$		.		y�xgR����Z4ddC;)43)?k�nB.Wv���\?WCxyeR^��xU�IR)/Ud��٪�{N(8t�vtt{G/ARAR��RR�Ö.B����Ƶ�jj�\@Q?���Ɯ��͛�j\\$\��w��ͧ�����ٜ�j! % 'ge�^<Ri���v�t%Et�MtkhvbBQ�����@2@++!@\\QQ."8EZd.	yWf���g#/g��a:'7FUR/#3r�NS-M����[	U�RUx<)x��sZUUUU<:�{���];R:R��U
			#RR^�sr����hb�՜�՜�����wnk;Zr��������ƅbN��������~����ƛ�j@$ 7<) ^xxgRI^��x�iH$	+}�j+66\}jj����}�\Q@6}��w\+6.NZESSd..%xϾ��eRI##:e��aFxg<<<#Ky�GG-J���� 4Xe�x<)4G��~�U'<RiAasx��sR')<AUU4
A^^RRe���H.9��յ���������WXif�������Ɲ�jQ62W�������\t���������j@.+;da%'Ag�xgR<x{PC6@}�����}j����}w�}\H@B+BH���j@6	.XSSE8P	&4)<e���yUg^<##^��uKRIAI#<eyKyZNNbvJ
PexxX<�����G-<P RLGd~���sK%iX;#R^^Ae�vH\��Ɯ������Ƶ~GPkm������Əjwn\B+[������wn`t���v}����b&-id��iC'3gx^ugRKR84$\jjj������jwj�Ƶj\jj@@j�j\v����@9@+E8EF%			K3g���{oKxxA#g��a:##:KCU�d?$?8)P�e43���Xi4);<' F�rEi���a^< 8"CdN7)'3)

^�:3Pi8 Jn��՛���ڜj��Ɲt~mt����Ɯ�j\���W2[�����wj\w~n~Wj���ՏQP���xa<)3''')<���x�g3R<?;2t�����ƾ�����jj��ƛQj��j��͎wjw��j666!%F 	)44����a<UxARp^'//Aa::FdG"%?dx�#4��F7C7?PJ7Gd������^KK<R)%&WM28t[?)(<a^'/��EiE0��Ƽ�����������ï~f��ç���jj���+!!k�����jvjjjQWv��Տ��?)Ux���eR//IRA##^��x�gK)ZXtb��վ���վ��}��j��վ�}\����հ�w\jjj@!+ 	- )G����K<'gx':<^:/#^ug'33
0J;����#RiiCCixidi�����ß�eKK]<2�vM?f�i;PCUR'U�7)EW`��ƛ����������ƽ�id������}j���jbt�����nnb�bj�٧���i?4R���xyxx�UK#:e�xx���Ud������;��njn@n�nQ��ƾ��}j�������hjnH.		%	$2,88idE���a3K<<47:/Ay�:4P)	N�N���e'#Uo�{e�ii��«���л��')3(%2hvh2bv��igUed%k�ҵ�����������-7]~����jj}�Ƶj2n���Ɩj\BQj�������v-%'3R^��xgx��g:#Regx��������������@.&B@6nw\9j�������}�������wh66+!
8?%$;8?%0i��-;PG<GdiG U�ei��d$ik�i�gR)33'ye��ga]e��{���Úii)C[WtwW.+jW�yix<%�x()9$v�Տ���Ƶ�����مjM)P�����j���՛j&@vw��հj@6Bj��wh���N	g�gIKuu:R^��uAUxooU�xg�x`f��jjnjj\@+6@+Q\\Wvhv�\��j�j������}\@@@@2 -8% %%8W8Wf�`G2NFCPS,&xeC)7v����tii�ig:3):3UxeeRaU3R^e���{d���P4)<)4Ut��jQ2w�$;aLZR))XrX0J[2b�͵}���������ڰn9Cr�����پ���}@+!\vw�ƾ�\@@W}}}n����%<��^IAAIK^e�xux��x�aKR<?eH[j�j6!6H@@666@Bh\BHtjnh���������}}j\Q++% 	
$4;07 ()"%9vM�t`9`S�� 8[J&	..H.
CdUC)3X�����rX��kU]gK#/R<3<RgRL3x��eUe���()iSk�nb���k
CU3	
	 eG-7P9N�зwj���������ƔN	%tt������՜��\6\t��ƏnQ@jwv�}����k?G���IA#R��xxKI��d�d47C-?tt\hj\6@@@@@\9.bhHbbjQQ����hn}jjj}��B!-);4CC7))
 88i�Q�fMNNS�[[8kh?62.		
Pd:(N��v���N�x�rxxK:Ax����x:��ԇax{�xyCyd[?Bn���?Pd:

	
Cx)) J��wnj�������о��N%S�~������ƾ��\@.hvh��jQ@Qjwj��}�w�vt�ýe#//#I���A#A�gadGSyiCPt�w}j@Q@@+hwj\\\Q\hWt\bQ8wƅ\hQjjj���}�\+ 7-CC[X))) 02Wkf�f9WbfM8$Bvb)7'i�����dSiXi�x�:#<R������U���eex��4KP)4t�M9M���t S;0 				)x�)9��w\w�����հ����Z	`��ϝ�����ƾ}�}Q2bhvj�\6QjjQhw�������~�i/#:R</gs�A3G:i�~~��QHj��j\QjQQj����jwjnbBnQ9HHw��MWj��jw��j\+&
)4;`idX)))( 8F2bbb2Mbbb992	)))XtttH%E�����<:/I�������x<g���Ra8 4Z��kWh�vff)88 299?8 	:Z�<b�������;��nj��f%k����}����վ@\�w6W�v���jQQ}b6b���jv����Z'<Kx�g/##^K:a<Kd�kf��}�}�}n6j\jj}}���jj}�n.HW?HMWwnbWv�������\)4)XNJG74)%.29JBB2?B�$&2H..&%44R3<ZriC)"8����G''AA^:<���xeLAes��4)?%8NG[~bv�wt�i:.++H6\@ktt[2 )ZiRF����Ƶ��Ə�w2b��8
`v���}j���ڜ!Q}hvn�����jjj}jt��}@Wv���[7)g��^):RxsJdt[2+�����wj�Qvjj}}}}}}�j\}j2Hnh[WHWkv��������}@	
7<GJXCa;3 .?H&+n.2t8%%		
KR'4x�G7E?��ti;)F)'AK^xXe�xU:<eyg<3:8%7~dEft�vMPGCC,%$?w\W&.�t-)��A<��v��w��w���nQw�~	Cv����}�����j@bM�n�����wj\��w��v@b�iN�N)'x�R/3x��y��b$&��j��j\�������}\\j�}h@Q29bbWH9.B������}��Q	)PPPXtWP<8)
		822$WW	 28W'G()��d[v����i%):I#xsx3I�{i�fb{LR�G<7PdC��N?t�w&&..0H\\2";)Px�:
;b�H�w}��wj���bk�&j����՜���ٛH	B)"N~vbv�BHE��w���@@��b?J;%7XX)P����ٵj!j����WN��~NEvtb�\j66B6@HQQH9?8Wt~9��}��j		3GCJitv~kZP)	
	?v?2$0&		7PK(3-������if? ;':��o3)x��r����K^<ZCUZiS[MFv���.	2.HHBbjQB)(3U�U/)N��?2\�w�����v$;k22\����ٵ����ُ ,NNbQQt92W�����j+\��tS?J;;P;^�Կ�ٝ}j@6��jW2$.9QHj6!\j6@QB.?9bW?���wj		4]irtvv��dEZ)		J?...	
	NJ-P7 �iJ2`X80%  4(:xxR)<o��X���<K�ie[MWJJJ��ht0(?t���vwB+;?GPUXC�{kkB?���َw}�[2W�t��Ƶ�՜���յ�\%SbNbb@`$2����ͧ@&MtdS7)G<Z<;)R��̟íQMH��ͰQ						29n\6!\\+69B&8!92Wt��n	
)ddf���b��ZGZ"%"2..!&%2 %E0--?;);-~J"%88P;7'K:RRK:i�i�Z43<aNC8 F[bv���i)e����bQ92$0?[be<'<3��`M0H����nw�w[EW�����Ƶ����Ҿj2.	,dvf`nb9%?�����n66Q?077<GCi4Rg3<x���kft9@@�Əj+			Q\nj�6@\6.@+!&&!2bWWQ
 E~[f��b\wtN`?$$%0	%"02!@6.2BM%;[9f[88-)-?�i? &2NN[~�Z/#/��KR�U)<'))%%?��w���Z'aIUrrt?.262&8[N�[P()
JrkJH2H��~Mkw��t P�����;��վ��8bbBQ��&8Hj���j6$..2?PCeiee<gARKxG)FCStN\Hj\!		N�����whj.6@!!62+6BQWB2	8Nbvtwv\fvtbfv�M.%$?JH@.&MwBb8%8MJWtt��8$%).G{kW8F[�tk���xA'KIAx�<'q�e:�<)),E2HvbtH[N;P�^g��N,$%$[�ti;))))GSEM8&Q�b98WH?X%X��׻�ư���B?H%
NfH9��Q!Hb����+22&&$bti�xxgKRKR)::-4C~�fQQ@!						t�����jQ\Q!Q&&H8HQQ@BHH&

%f���v�vftWbWv��b0$2%M2?Bbh�[7
)4CGEHh~��tJ0??Pik,,?fdfk���yxa3^^Ko��y��¶C/�:Ue)P[[FfMJJXNG�xA��X 	$N��PC%;%N0JGi2&W@;-EW)PPi�����Öt.%	
%7)fmbn��6n����j!BH22.?���x<:7<K<(KP4,���\v!++!			v���B.Q@j6@+@B@BQ\B6	J����nvftb`bn��wvG$&.?2B&	[��[G)ZZ"E,W���d?BM?NN8,ZN{�iirC;XPe�e#x���s����g)i-)4)e��N<8m��dZ[<U�G)
H��i.- ))N; .B8
 E�i)Cids{�����W2	(4?7kv����Bn����j+@BB2HWJXii;g<R<333')�̰w9@+!	tbWMQn\$MWMHW@B@2		?w�����nfbQMbj�ww�W$&%2N??�Nt�?)CiF,F9t�Wft22?PNG~�����fCZ�x��R/��3Kx����R:<gU/)P��K37N�ׄ88Z7diRHh�[; 7;%.,GF;CRR<3F���[	)LXfbtn�jQv����j\\6@@QB$?%)UX3'ReK'P����wj		J8$9.0.HW?2WtfW[H6@!8t�پ���hWQ9btjh���\2&%J?b[ ?t; K�d-)8k��tddd;XiPPr��yr�yi��x�Z::dRFryr��xR3<RPC C��^C��Ѐ0M?;C)8���N.%4)G%&&)C^,H	4-Kit�vn�������wj��B&.	PL7��^K����H		0HMW ,9"FWf??8%0b��յ�}wjb?Wnv\\nwHhW2J8 $ ; --[;:{iJ% i���fEdJX[�eZdC:)7]ddr7eRx�ܽ�xeeeAPCC?()R�^::x�Ϸn?J2	
,F`tJ?[8Pi)4id;)
 4Z3);Cr�tf��bB����vjՉ9&%)8Py�ZU'4itb\&		;%2BM? 2CZ[kikN[H%"����j�w\jwnWnHv�nH\2nn9MB$	):ggxC,FNS7��e<CRG;Zi�S))<N{EC�k����[Ce�eXPGy[PXLK^<������v9
 JH89BJ�P%i�K':x�i

-3^3/gd%%!6&	JXFCLqiGf�b.�����h\B	Mv�b`F��x<R'),WvH0%0EEJ8 d�������̢:4t����@H@h��MnW.h��wj!B\QQJ8-dx�xx<-)<,Giri�ϯR^R<C<<��q(RxU)ZNi)CxiF[���;UxN0NixxZ4I<d������v?,%%-);i���n���k0 aee )CCKdxR����������j&X�x7)CC0.EkW9$����h9
J��t8;��tC'^<'#:C��n		-`FW������iGe��x')0$�����b6n���n2WwWBQ��w.6WM[f,%PX<^R'3;)-?������iARgR<<eZdx�y8Xd�dEX��i%t͔�h:?PXtPNX<e7Gt����W9?N9% :)X��כ�Ұ�b%:Z'

4e��y����sr�����\&t�S'-W.E�ttd9$ % q