�
 ��jb*�nZA���8��{�������r��-{ $��
*4�,A�Ck�y�V��pY� �sM�Zp�i��++S�?gF�E��,���E�w�q��l�|�{����%�+��E��kuy.,��Mg�'��k�jۀ�ӊ��"�.����6�����k��l2�e.����q��¦b���ާ��Fq�J͒���r��P5�Vs����dl�K��}�L�:�U�dt⍳���P@��0��Nÿ�t�U���e�f�Y�ږ�hr�s���=V�U�δ㦖�B��]�}�]G��8ǎ�6n��6���t�1(@�V�Hd>�9#�����X��}����+Q��"���ŧ*�����;�{�R��|U���OH�I��T�i:`)�9yrY����;�t��J�GG���m�I�4Tc��p9���|���GǌF����8b����tP�BS�;(�5ⲝ��w�4���QL�Zl`Ƴ�������E�7u�ZA7<�.� [��5�`��J^�v����u[ty���؂,��kE�$����z�t��eZ�.�R�����)߂dJ������gzҿ	*�1Zdbt�m��x�2sNnd�*����1ۀ1ۀ1-d:����~��or�MJ��3��(-�����3sl���!�,���,��v�?�,-#����`�ϒ�g��U�,,{�\����Q��D��6�+g7���rn�P��`S�U��*�n�n"�I,�.�v��'n7hi�mw��	��g�e��V��C�p#��TL��p�V�����ec��
�����I�[4���ϒ(ѿ�dz��3��-5�� ȭ�)v�ǼL��t6"���ؾ�n�so��ƻ=�a[a���b��#|Z"5��A~�Ɉ����LN��O����
U���;[=��g9��
�I�j���;���x)��2rM-��P�n�!q�+g�9�)�b^wc+Ʈq�$�4�=�n3�un��g�&�n�h<L,~@�l�@��֧`�o��E�$�����(>�Nt��'A^���1���&�����Y�)��<dnŦ�c���f�Xp�U��W�������8����c�!G� ����l#�dϐOio�� �Y�Sñ:�qwoJ�nGL�@��H-�o�uLN#����0���J�H�R���J�iT��2 D6�"������!�vPA�YG�I1�/�5�Թ�s����nύe�}jfȬm!�UI��ܸ�c�L:��'	��N�I05���]9�������g��+�JG��dq�F͗�uĞ$I�qJA�y&"p�W��� ~��Ol��\�	7KM���@l�<�B�鸰hr�� I�\��/ґ�wQ�q����5C�o��O;��	�'^?�*$��q�*��܊�L6���'
��	e �d7C����n	�����;�=��_b��8)�Le�'	����w; �|�TJ�����o\b0� \u��M�L��:�_s��m ���a���Y�n4�
[��mZ�ZY�E�a
.f�z���z�"��C�����<����tܛN_���d`����7��ʿ2tm�$�w�:���e�R�UZ
<��:UN�=�:	  `č4Ư&@.� q�㓬~�Ƶ/}�)Y7�+ ��}��$y����G݇�+���*��A�[%s�}n�k��o��-V����;2���9�Ϳ�G#.�j�w�C2��ӑF��9<D�h�p6�<]��P%60�vs L�/�xo��F�E��������O6��[n���_JF};��?_��_C�D�)���.�n1�7���f�����eB�,���G=�>d���."���c"϶��O5����1w%z��1��tu��".Rv�s�z ��p��J8�ihwE��g���͞H�ٳ���T��Z=@:p9�3�A��^��IQ���d����P�w� ��(ڂ��V;�yZN�Έr���8QSɴh�u�����������]F������[�	�9}���3�_�Q�&�_f�4��g�gn��P��������\�\�<�¯M~]��G����W�y�m�A��v��ѽ�L�¾���v�7������x�C;��2�����L�~�T�����ʓ�(�2����c���qo��-��E�D�Xǲ����F�~K3������	z;�{����*W���"���ֳ9a`�o"��������ĀUHO�����)��٪�ߒ�){|Ɣ�C|zH�f�}T�KKO�a��p+06�񚰶���������������5��������dO���ڣ�c�/�Y|����b
����j�&-����S�> �9fJ�2W���k	��{0:��oS�L����!�����bQg�s���q�� p��k=U���-�"���J%ҏ�Вn���a9gJ���~k�����}B,:��/Or���x��<�뷺�������K'��f�9ޤi��G����O��л�u���˯�.��+���O\��p�T£�3��b�H x��%��� ���G��2��
Rĥ}�4�@:Sä����ᆄ�5楅m��/Säi�3�ri���%��nu f��������f���1\S��JR��`������՚p�g�������I���@�P�v����a�s�n������2��%yU�2'd�a%���ԃj���F���'z�6�c�b���}��n�pn��Z��K1+��wo���b>-Q��ۢg��sc���Iu'j%�6�U����}�I��j�J$e���O���Q䑳�uI*ʹ��H��~��v*�����W�e0gNd�AlU,&� `S�[�\�������$T�-Q����	1����\a�N_�.^� y~Ae��A�N�_z��G���	��Z���v24�g�%��`��0��_dneo���G��	ej�9Wd*i��y�^O,Բ��N��N+���D`!牫0����ks�'"D�Uk�!�����Ү3E��Z��a"{��n��é<��1L
Ƈ��;�fɞx��\4]g�$� �l;�ȸ�����w3�o�g�v�z�D��+�	8�*��p����$��6
�VC�ӌ���t�`�Y�up�a�^��[����i՛���W���\��|\=�c=|oB~Y,r���z�?�"^��i�k�9���Q�v��ǇQ�O��o,��T�}{�Ͳ&�4hn�e3�x.���n�{�'}-���!w�H⯼�d�^܂��#��k �_��/X �o7���.6�Q�����&^��<���P���[��-�<��m�Vq:�Xm̻ә�"��׼=��ˤ�z�\gH�(Z��c6
7hͻ�X��yo��'��sj����^u���}��FVa������٣A�<n,^�$f�Z��G;f|����#�l�oo�����;k����3�����G��D�h��Hl�3#t΁ǧ�b�����^z4��𝄩�k�ԩ$�(A'v}�d���T�k톯k\�Az5����h�C���umJP(�G��y�\�G'��,���E�����;��]���b����1��0�k+�\�(�}����O�������K$��"5�'e�S�Zg� �h��Ԅ��N4��Ǎ��S���`�hg�҇�p�!�µ��ƪ����n.�

0���V��tz��oD�$#@��W�H�pƷO�rR��A?_���rt�3��i��x�AԄ���������Q�m�/����p�wk�G'1^R�!����P��,nG!��(`�5��'�����T*�T�o��w�"���ǉefS������D�m�oȂ�4�"�!�߻kh�����sӂnb3B��:!��z:�Y�=L��a�H=15��QL�f0��l�
��"i�a���*�����&efǢ��ľ$o���"�^����%h��X���O`����T����$��d��5<��Vc ��1�M�`��n'�UL�lD��e��we�Yl<@н��t�W[�+�w ݘ[f\7�����+K����Q�0V��c�JC�N���z�=Z�y,A��<�<���ZW?��|�t8* �Z,����y��h�[�d���H��y�2��{��C~8�f-oOQ5W�{u���Sp�EE�=\d��R,-D$�0�՞�����~:�I�UeO����_l��Зy�N!x����v��0�8g.͂����Q��M����I����8&��K`�LQ0�Y�B�ymɌ�B�>ĩ�I��L�����U+��}���%[����Bu?�QM#aҚ<� �S8Z�J�s�s�-�Tm_�6[ѨI�ݑ;��Y�����w*����_��I�,4 ��ۻ���E�X�y�.�|�$�_-%��YVK��a}[�C����m�*�: �e�?�vx�_�/3�˲��/B�1��<�!���v3�w�nJ�&
�?.[���-��~�x)CiU\J+ԁ��mC��p�?�+��ZK6'G@�ś+��0���V��OR�EN*e*Og�w
r��dz=��K��[����V~���0,�u�o��^�0hp�d�U���BB/}��9���e�<��ܑSm!�����j�_[��5�dD�f��FSA<%��w�9l�ϖR�o_f��Q�S�����IT��@ټ��|�Rʚ�d��ѯe�9 �&Zf�I�0F�sݿ7���'y9�9���'<�,1��zۖU��sP�L�[�Eib�d����u,!Z���'�'�c�ߧb�f������S�T��b$c�gx��C�csQ��x�gru��+� �o� ��w���v��la����F*����n����C��8 B��$���$�|�/%��cg��)��@+���(��K� B)�#eS��jR�`��4��nu{'0��^�`gǌ�l��]�U�	����H<�`�1aa��tRP��0�Tھ�	
Q���4������T�^�4b�	���fG��|��8�V_?�������ٱt{V�&�̒L�a��rX�.>@��_>B��,C+����_��9@�K��-x��+{�K�]![-Ǵ��}�|���-���Aԁ�,t�:_'�V�������.��1�֟ǂ[)H�'V3q�;�IG4�&�T��s��^�`�-(�˷����du>JR��
	�,�h�V��L��Cm/�B�p���}�I_�ў���jp��?��3��t"���S֍с��ɫ'.{���|�����p�׎�w��n�OS�7
3��5%[�� �B���%?h`���lTL�1G�7n+To%�)���s��`��0=a������j����ʦ�Dt��3��ޑ�)�H���1�j�z�*)���V�W8�q~k����x$P ���ʇ�*Tw��m'-��X3qK���#�p� t߁xa<�i�vF��M��$n��#0E�G!����W�½���	Z���Z�Ci����ݱ;�O\�۫�Z���L�Ã�K�㋔N2�� �����д(�z�z���AYHg�.]D���p��P�c��n]$��bQQbkw�[�N�*�ŵ����v�4�*�'f����ƙ9,��%g��9iL�.3tٷ��W�0�� ����w�_�D�w�k*ف��׸x�h��֠��v��N؏�g�ɀd��3�H�e�{n���)�7�����Q�P ��%�5/U�Y݋i�"� �����c�v+��=�JڒP���S�������S&�Wh������M7j-�q������4�a��'��8Z�6��f�e�N�
j-�Qn	zK@����b+Qi��z!��4}S������L���|'��2�9W��%�J��@ݑ���-�f���5�Nl3�z�OT��2�f{���j����|'�.��i��G[�W�[*������A���4H	"�"�Q&ӵ����`��H�Y�A��@"��f�I8���HU����m��!��J���
�e���Og���!\��8�D��	#&���`�4��x���O�<��.�)�b!,Q��
�e0�ʁ?^v^���@�O#Dڐ� FPh�����N�Dۗ�'y��� ��z�IA�(�R�l�CuC��W�H��
�e�(�Id����$�O��} �Cy6�-�iFE�g��{&�d&ʉ������M�LZ-�����\-��M�E��}�HᘂQm�� ����'j��Y��0�gJ��g�\���&�l�U(*���*Γ�3��y+mz�G����zP�z�T�`:�	Jj�Q�C+ ��o!F�>�7i9�6n�� �pIR{kta1+�lf->��1o�[?�>Lt��\M�.�Q
y.G�t,M@�:�����z~-��9�1�@pA�Iȓ`-�#��{����J���Ҵ�y�h�^���Άl���-YN-K� �>�(��f�J4齙�f��X�5N(��HI��P���}mõ�R���~F���W���/���<.�2����!�V��Q�
�y]����p"T�P�[�{56y,φ��QPWMϦ�-��E�ʧ���67�j�@U'WRv&5�����V�qp�h�����$����_��>�y-���u�e�ΐ�5�����{��R��t��o�P��atĢl�'^F6.���k�T�eN�����zA�}�Wp�'�ާto� �jr��@�>��6�B���'`��z�&&��Gp���wjgp$,�4�`�`�̑�}t�M���z�9^*K�ġ^�Ɵ�I�i&4�ЫR�R*�č�N:eU�;�4��|&����[�h��R
��>G�Z�Yi�eA~ ���A�qH*	�R��y�1V�s,���hÔ�}�#����ƾNl�9i Y�9�~��E�k��0��׹!��d�c��xtZ ����O��40��Id�8˗�\�t��U�j1�l �«j.��A����?������T&�����&a|���7$d)-�N�?��!o,d|��"{p�H-w|1��A���"�k� ���E����N�D�(5f�%&��rmѥ��`�k�� dK�ׄ�""�q��#eQ�SFm,d�с-
��\*{�,����Q cS�ԉ���``$������$r�L���Ǟ�[��ؕ��D���U[�Q44����E�&���W��]�e=�#�3�!��_�H�m�+�V^����aT���K��s^3G�}���d/��FqHk�ڗ���G-J>�S@��~��\���T���������$|ǥ ogJ ( 	Әh���n�6A����l��W�.b.��!����PƏ�V] Q��s���b��j�Tw�P��/��~P��R#�]F�5��E�v� ����,�ʯ3D�>6FO�Zь�9���@֑* ��m�l0�k9&�N����K��5M#�%��?��Hס��I��)O`���>_uLa]F;�����P]��O�:���P��Kف�痚5�nI-�G����7T�)zFq0]�ḿ�Óc�\�^bs"Z"�˦;�/h)�n��te;R��P�����<�H��"g�;s]�ŭ�W��.�\��+)�wL�x�b2�	�Q�,4l������1����@3�5Di};s�g�s��h�����ނ��q�Y��Z���ұ�f�c!��~�k�1�TSU��.�ԉ��.�XM�ip��K���y#�R��}U�Eb�����*g� �b"z�C�����C���Z�z �j��Js]�}!?t��݃�-f��f���s��q���^I����ﬥ�A�� �!��b�'����d$j�Q�]-$�&h��X�7�e$�M��� ��r��ce���a���Z���#��r��rMMJKom�J�M,x��E}J�}v���G+G��M0@�,v}���[�^N3۟3�rh�$��w�T���W��nd�E��GQ^ ~[�rp+O_P�Н��9Yub�%,֌pm��K�*۝iB�GT�Vʥuu8#l: �3�VJi�%�V�U',8�S�(�Q�P*�
��Z-��9��{��Ez���C��M�����Ĩ��tؾD���Z����J�VlXN*XcP!�4)=�1�V~h��X�ړ}.�?>��?>R�j��7�Ȉ�M�8����ѝE�$q�m	�Q�f��l��75�y���"����kh"'�&���M�e!�X�7~/ /�
.�</�$��@�P��CC����E%���� �����"{#h���j�A��h����-��p�X(�hc)����������~�R�1c�6�hJ؅��&�4�m�F!�">�-�#g�
��h��m���i�s
Y�/("SJ�b�U�t�l�mW��B������U�'i!.c�x�N���N�¸y�����W��O�;�/��L��A�dD{��.jecG�Ta(�_�z�`f���;� �������'�2���-����5�|�'�0���vt9�F�p6��u��˖�Gv>�	?�H��O��5bƫ65^^`�|��u��း�=ߌD½��'��ƪ�N�䞄�3��Ɣ�z��6�q�k�lf�^U�-|�ox##T���_�ECI�K��$�0;�S��O%�"�TB��	/����9�F`�Y�A[���7��O��:�b�6��(�}e���Ww�����)���J��M�v��H��t�4��n&�諿_v�����`�i�Լ�̩�a`��%�ku7-<��;�ʶ~�M�e\����O�Ƌii7�n6��)��(���cz�D|�%~�%!�:����$�`]��@���G������7�X]����(�{�6j�&_�
���{jEwl�F�,˕R�jiǶ�e�KM����1�w ���(�s*�u�K�c�b/9�s�w��2*H�)���L㵎g��=��n<	]O��K�n��K����45l�>9�P�y�6ZK1[p��U��`%�������'�D߷�m���̇a����������b��<���)Z\��C��굠��h�e���L��8��}}������d����5�e�7���\���d}O���b"�g�TJ�`��V���(&m� m���
D���8�l�������5�������@�'N>'�3�%��P�4�z��q�!d�=��q��_ !��}��N7��a�Àj2}>���+q�%'D0���o���om��o�3͹4s)���Xe��\��wfK}Z�A7�ˠ?$4���:��8YV��y�(u��}yw&&岑}�q&���WԖHb�n�=�#,L[i�hl�ʶU~��E��	z�Ţ�B]�-�l`�y�����i�φg�dέ�a�@�עj��a>�tx����%����%ܓ�ō�k�/�3���D!eT���gA�8�T�@r�/ i��} �D�G1�y�����.0���H�DAF����:cd{�V�bC��h��ߙ�spGh�{XƬ|c4��YI�.�0{h����������n�H�g7�Umd�˔i��m+H2-XvLh`s"׃�}�^�D=��y?����wV�&���Jz������f����v�Cڳ�N��m�,�:po�tr���M9I�@��#������N 	���杌�J59Ƣ�� !�����|�T�枓&ԍ����Y�sЕ;i ��'s�NaR�%Ϲ��.D-f��t��o���h�8R���u&y6+݇VBI����X�|��ӯc��4�����e)�tC��r��@.��ӤH}����j~æ��i(�v7>�8�r���#l���Ҥ�Z�E���O'�S��C?�Q�Jk�M�pC��$<��"�=��e�P��3/�>"t>����;�3���Z���+�U��V!@&��ހ��^�ǣA֧nIb�ߴD���f�@��g�����9
#�A̖.c]�K�W�W���4�Q`�I���"�E �J�𒝵�+�g9}�V!.�7��$B��e��	s��0��)g9�d���-u�6�VS�M9�z���M5�Ot'���°�H�%�O��lΜɌ�z�*!�}��n�nٸ�m��#�m$b"�@̋{c�|�"���orT��I%��GlgWa^�'��9�?2 �P����U#<�xFe���ƚb���Vf�KU��� ���J6
�:[Ϛ������`���ɠ�w`�������q���ԀN�����F(|��ڗ�(뱀�)P�=����(�I����[���=-�E��C��`RBi0�r����n�8�#7N�	Ϯk��j;�`���1Q�I�6=-y�&t�E�I�	�ݍ@��V蹿����E'A���f�Kж23*��@�J�P��h���Q��@4�z��0���� )Q��?�Q�=����_\Ŗ��EU�V�o0H�OɨFOx=�h�C�sd��`�O�.�Ⱥ�o��\������(yT0l�eN����ԇ�p��
��v�t=E��1K)�[|��uɾ�0�3	�)�)Q�Uo��9 ��;˂��v��b|��֝F~f/D�'�����0(��1t�ykh��Q��9#�?�{�[��8)�\��+ܡf���Gq�,��8�F��ygy�Fg��X�$;��k�kj9�?�Cm8ޘ,�ŝygmy*b͎����E�V�!ճ"qjb:��b�!r��m��`���#��}��Ra�������h��`�������=������,��j�}��&��@��X��iA�5��G|�o��[u�,�E���(Z�b�[���dl�Fc�l
G�!cʗJzM3@�}4�h�ݓظ��\Y�P���d<2�� B���cB�c:&l-c����<\�Q�l3h�{+ee��p��.C�B�l�=��������ŋ�)\!s�l��ڂ��I2���kXq�9�m��<T-�yۋ%3��y����v-R/�$[@�����;�b����Q�.t��}�j�G�g������Pѡ���M%l�P�I���g����p��V��@Awݻ��}�DF�ǳ�7C�J�0�YpΙ�E��"�p��p�:��ټ@�ZlmzTS�=�=|��B��-���<�}�~�E������M
��� U�4<"2<l�c��Ha�6gENn?ˇ6s��M/.!��E�/�"����ԏjV5���pNn�m��;�J؆5.�H�Y�p��$��%��j�Uh�9�r`%IՆ���e���X��@���`��Piv;����k�o��&��:�%_�$�'�]�݄
!��&�4�<i��6��62��"Q��F��;׭��-}�Oe���gg���ƈ�y�n�3��PY��h!F�;z�痺t��eJ|��T���k�$L>��-!�7ү�����h���cy�ˌ�� ���<��*���d`���&��m�hB0�HFhȃ.��<��Ь񳿄+��t���g_�3M`��lSb>c��Y��x7N�AP���]�^�OM��H�Ow�P�y�^<h:�����"���D��ʿ	F�E� b���u�2.y/�%m���iw6�r�A_�DRCei�sT�r|���Z�r�1J��0ɦך(X��U]�W ל���V��IT	&�N��w�wU��.�s�sd+�ߝ���*[�r��&S(��4`��P���N�������w��4�\���쵄�=Bp�������"Dp��;��ǣ���{�5��>Y��B*R��x���u/yս�$ ��T�Ϋ 2Jy��~�	K�K)V8f�N���L)�~/�(A�ә�ΨL*Dm;��(6���?�f���/z�T��u���dЁ�L���5�̺jH�S�����o�û���^����My�Q����1�� �nWY#�,h��8��<8�)�T���ݐU�W��	t�(��G�������ˏ��X��d����l�F*U_�뺈�{H@B�-�{�BK>�ڊͼ�-a@�au�hh�l�D*IQ{�\N���~M5�=����S��(0t�u�U&m���>{��6�����x̷	Y8ړ��R|�{w���Y�r�B	7��r�k9�˩�c)�y����r)�R�����ᰊV������c��΅�������ֻ���a�}���n�c���MrU\� ��i���N��1n�%ea�zV�˴�rw�sN�4L޵���t�)J���bz%K���#�ʻHSӛ�!ҦE��u�/���~������ ��=��;��:h������aogs�(f�����ƾJ�5�nt�a�ΰ0�ғ�Jf�G-�: \��3z�y��4���G)ӌ��A'z�{�����񨲽k�p�����4�HO����FzQ#U�\f�
r��8�O�9V��6�<�$��}�����p����<��<c<�T�{Ib�����7�(�:�oO�j����:�7���Ƙ(:��b'�j�w}�(�����l�h�����؇��f|{�½��'��x�A������%?��:�D���Q�.j�����[��\�	}e��@�H�}d���	�.[�;�O88�jȉ-U*-�p%2|5n������a[&�+8Ԇ_��T)u�:=jӅ��ŀ���f�W�NOY�7�RjwVP���E{����iu̴������)���K0u/�B�~Ǌ���191�W�wL,CާXe���G-$���S&R�q���b���-��O�V��c��!��Zc,�
�H������߂�@W���VtM���ȇ�@֮<`�&%�F�����-��~��,\���\���JF0a/�3[���K��g&�ۺ#���A�'7��_�,�=�K
JB�#�:r-�R� �@�h8�̯D���l���Y�����%vx�H,TMi$��_U�)�K����s���fZ� ���]r�kMп'J?ƥ7Ļ�Ǻ�4z��py���mH�\Iu-m ��;!���4�c��`��?7���.�g��D��-Q�f��e�Ff���V)�l
.��;(�v�Yp���X��2y;���;�;]2���!�Q�AC<ߢ�#�xx+ �i�����o��������h���l:	ТS���C8��.f���d�W&G�������3y+��"o�ǆ�uσ�y3�����9�/�T�SE�C�_�2	�f��%)
H��XY�k�j[�Jף{]�'Be�����xB2A7�)�M({�ﱈ�͞���������5`$�U�6A7\�0�N�@z�S��B�Fj��9=����?s��R5��S��=)�"�ʙ�A
�w0�@l�S��X��B����,`�f�%`�d�Ӽ�'!Ax�Z�uE�yL����ZZ\����v0�L��ϭ�j�\Z���'�U�_
t�U���
��¾+���<�i
*<c���$��=bN>k�k7�	�u<�Y��:Nua8!a��u�Y�!�X�u��e�&f�B��b�J�Mgb�zwbӘ5�aԄ.����7���g`�C��t����7�B���a�����ZM����v��$ct���kw�Z��!��=ӞƛB;��_1^8��>R�hs�Z?.�7 �a���Fs"���@���<�G6��&��-�%����#T\ϊ�zpܽV$�2�+�y0Z�!��R$]?�����k�����W�[U@�+�!�E��u� x�P�����,&�E٪�t�FB)�tY��Qj�8?U�F�ȴ�]�Vɜ����z���.)��@&��?6���m�6�>��T)��2��a���(*ED��z�Xu�j�8Bo@3��K8mnk��x���q��]#z��\��q�,9�l�G�Ql�aF4��ʚǢ��]n�͒g��&#�̾���%���%�����#��^��PQ޼/��fq��8a���;�Yߗ���9����L�`�v�l�V��`�Jre�PP��tQ[S=���k��,�mC��m�J�纟���@c����n~T��	�:����t[��>��X q���C5s=m�t��S�
��<�� U�5�
����C9YTQ�'4�~�%H�"I�#N�$O��;\�}T�|��-��Z}o�·�	����3%7}�����d~[x���/�b�����+�lFGԥ�b��W4˶��Q��/R�u�'�x���1惺�{��x�5���[��ǟ�w���ߛ�"�W��
M�sg{��(*��b;���}�u��$en�;cq��O��c*��;̬ <��ڻ**����;�l�X�'�b��?�d&R������ߠ��M�{�aإY�&�g6g�CҚg�Me�ӛf� ����Q�b��5�'�s����M��
3�0�Q�$����z�s�#�T	S�@���Rs���"����T��ܪQmɑ�o��f����JgQ1T�`K�͘��޼c���	l����0W=���!��:.R�n����(����,�HCW�6�U���jXN�J{��#�á�P�]�@�?��&��n&��ÿ��.WsQY��g/_lY�T �P$�N�ei�6g�48C�~6�'IRjg~@��Su��ssg��օ7U�$z�Tj^7f*8㼙�l�*��xrFl����_��\��ZM?;�5}H���R[���Z�;�?2�Y��� '*=�Ơ��2��d5�C�Hg�1�Bu�(�`�fģ���#�bģ�h�������:3<[���&`���K��Z��D��~� B����m��h�#���>������d�����r�F���˖����kdcDy�R�@P�r�r�Y<�Ar��Z���#��A��Ԩpg���n+�OH�Q���>��#_w(�����Gb!R/��5���	yE �6$�$�oErXe^���(���kIP��o#�c~�e��E%�ԁ#�}>K���j�-��k@�D��U�A�+�dU��H��z����u�" i�)H%��%�K2pb�咇�N�k�ݙ��T�����c�y$C+��u|�ѫ�2��B%n6M�]��lM�����J%���/�t.�zORq��p�B*1;��i�7xu+Ẃ����o�����*�g�^ႶlMzU�b���ng8�DQ1�A����l)�
�����#Qz�\��8����m�A ԰T�4���Q5��tE�\��1�0�o��:���	.�o�m���\)������Bs�g�rk�?��8x}���@�)�u<�E}"�k��>�7'�o�]Di�A��� �i�ILB8�b��d�{.rF���ke�] Nz-�N��a����3�Ro�f��Z8f��W�pKH˒q#_i�����<oqXv����4��_�:�{G1�o��V�A{`q���=h]�W-nT��I*O�Ӭg~�
=A�r Pᱼq����]}�y��5�I!Љۄ5X$��#��E�DT{�N�I�)�����f�Y�0���pR�%I)��`�a�]�����y�H���?D��k|G�
�����[�H�k��!����G�7�¤
��l�w`i2�����3�K�ݪ_)������̡Ub'�4"[CʭX�/-�h�ȶ��0a���,��os��?R�z�&�K`�v�q��Z�f[�1����h̴D�W���W��0��v�ˏ�n��.$9~��{�R��J�̫
0��^~�ֈ�[4�-�jgT�� "�Q ���!W�C)�w�F��3'�'5�}��|���_+FĮo���<9K��,��fϫO~���.�w������^�]�ǀU{,��Dr �'Y+�z/�]��˓z�o�A�k	��SmP_2t����>B�W���;DX��J���a�+ƶ���Zϰ9��η�AU�PY����:B�L6O+l�9��\0ML�ᖣo���j7Y��S�;Y�����թ��_�j�'%�ğ�~�
#�?B�%�&s�T��1,�[�{폗�Vr��''�;���SU9K���Z�sr()C�"�nOE	�:��K�W}0�Mj7j�u~�=}2� �Y��l�#�vw��9� �m�.�!�KG���=_v�@�;��(V��J���珃�}qF�@H�&�_u��������a�Sh��H�ǐ��tF3H���1��G�6�m7~{��t7~��"���5��}����?b�
��*6���X�с� ��j�����~4L� Ⱥ�Qk�~��a ����a���_�K	�p�DX�hT\�~��0Nq�^�I=�>e���j8i.ƲL`P;O|%�Qd�C�=炜���N���	,���V�$Ď�4j<=gM���w�×�q�0���@�N����G���h� L/�Z{���b#]�1v��`@��g�~�B�BC�������g!��������P����Bp�^�W��F�ʃ�@�yK��	~�idr��mg}z��r��i�N�Xʀ��ւ���,H��'��q	g���B�U���W.��)z���[R>��|B�`�VH�A��n`8GNǳ2�,�p[�#M��x=#S�Əd�����,��y�@�}ըG7L�Dl`�o��XAo����L+
�H�D+�L�&���N#�V�2Έ��F)���)����-s.�'��7���L��L� B���#�Q�M>x�x	R�M��
�e3-R���~lg-L)��|u��� ��7�t���ip��%Gv��J�`:Oű��۰]�S�r���7�0�<��;��p2
��x�,rV�:����S�jX�-_3�Ï��O��X�S�.���Ϫ��8C�|q4���ZT�Ǿ\L�pi�6$}����z=���F�(x�uZ���)IP��ƢO�|?o��A�>S�ޫ0�̸�����[Z����&=nVRھ�����oǲ��x�Z(�����8(I�_��5���N�w���&�?�苢�Ø�L�G;����h�p!�laׂ�0�A��N��� P|����^�nd+�A�@ٰV$$a��KA�!J�m(ԕ-��\H�<������N�����TS�������n�v,	�;&���N_���'���*�O2���/[��ʴ�iqN���w�����=n:���b�0��/.�$���Qr�����n�@������-��KXr�yA~���45�X��B�hڜ���]S�:�:�y�,�!O�k�M,�H��^�7v��l\�yѹ̀n��&��	�M8�;u�S9�͡���S���`5�[�V���kUwI��{]�6�h�n"��̤�ɂ�gI�*9��s.���\�j]v층pj���Q�Y�����>�%v^�����kD��Y��o�|ld�8��z^^s�@�����&����WS�T�et�Ԍ�=9������41Π?Zy��!��˲�W@XF����#,z�lG��k��`߀��N0���p%~�(���\6�Pw	�o�	4	]�1q�tD����Zg���i��cM���2���&x�+���}-y1�)��� ^�ξ�y�z����GƉ,�uQ���}������%���)��xiA���h�W���i'B9���)��!h�p,tk��h�3A���Wh̾?8&N���r���\�}u�~O�l�ViR&>�}��������
N�^�$�g8��ml�~�6_X�-��ی�Ku|������]x���EC��2`|���X���X��wS��T}Sp�m��3��'�˅�o�G�Yi;z�x!�t����|� ���.ƤC�����СiJD��G۽��������e��1Fl2p���d��i�2��WN������h�)'�-�hU{��2�(�%&ů��)��1�. �s��.�$�m����8t�ЄAg�X��e!E�Jg<��,�-��{�(�@��Q�Ⱦ��az�߄<��6���}���΂�H��|"��v4L>yO�,n�"in�����r�Ù�K
c��׵V�SŐ�ӭ�w5���[E}R��Y�4
�n̍��� ����u�M�� S�o�Fi�F��u.F�7�w�K˝�2�Qc��$�	˪� ~nm�D�Ϯ�fT���)�'��[�!0�IЄ ���{XG�XM��)�StQ�KNNx�`6��*�mL�_�v�7�|sN-U�M��YFM��|/����;��v#n��1a��'�\�0�F�e$�%x���?kq��U'�eh?�/�L�+��j��)��z?��w��`�s�aӔ��lΣ��f(	��<u����*��$��Zv35��l׍_���kg櫺�ʤi���p�8�)�v�Ð��Ifjj˽����QaA�J���6ނk1P�����H`�,XV�+~h<W"VJ�5�s�-o�:��Q#u5�q��wp;��v씬��I�s�󜲁�+:�ʙ�C���A?����춘;�;��c�hd
q�Ag�y;�Ag��>�q#K�8���V��-C0YQ�"`w~�����1�[�xR�oȪ`��hnս�r���a�
F*n��1�8A�S�E1�l!�BLu��M���?N#�� A���Ұ�N�q(�S+��]����S��`�~��%r���%���Ley��g"9f�;�B��#J��E?���~ 	��;J���Eߝ�B!*N��ᶮ�vS����pN:��q�qy��/��}�n=DS�a�S��{��l�a�؀f�%j�dӇg3dl` "f�����r�V���?w�n9��0�U� N�t���6j�2�٫�S��pV��c�e�Y�f?�*��B���+<o�j��0�w=jF1(�c����k��J�"�����pʻ��gЅ���`��nT���8�CZ���M$�gU���;F�Hkd֬�g�z\��;b�cc�&�yd����Fz�,�GCdڳ�w�U��ig���EW�;���b�\�b윪a�-��%r�u �u�������$�zy�e���V,���k�:��qGEES)���m�׶��ͩ�a���T�}�*ZK�S��F�]�2Z�%v�#ql���U��ЖI���m1��s`�[�����)$m�6� ������ڛ�>t�!mb3ד�s���DR⛒ns���;�h��m��*�k���M��׍�c�~�i$�y�ؔ�d�v�9���}��j�g�U����_�# J�R�k㟮�:�gf���/o��x��Ү�-wMWH�Q�����-��Y��LA������!��ϵ,$��:�_�E�2����кH8��>#�������qwf��8@�:�j�R��T��K�������7�h��Kү���gX�Y��K[�ҭ����` ���bP�r�[����'�PY��P�58���\��⥻d��&���i���� �r�n���(c�5ia[�bj9��s��ҫ���U��U�������o\ĠAbB2���/������j�������Y��I��}T�3��Ӥ�n�Yb�Ǚ���3�d�l��m:#�}k�e'Ѧ�d%�4��{ƞ�Ŗ��b��Aեe�j;د��N(��i5�uP�������Π}د�r)O�ϛ���N�5�� :�