���~vdX\`lnffhr���������hjtvfbjt~����f��ȊJX��h>>Xlrz������xr��������vtpjh|���rz���px�����r`VZbhn|���ztv��Ăbx��bV^x�l\h�ʴ����~xhfx���zhdvz���|j`jpxnv��vp����rt��~lj�����������tljfhlx�zztvzrhhjlnjrx������������pbbr���������|lfr��|lnv||rprrvvtx|xjddn��������|phhp~�������~~���~tv��r`XXbrvzz��|phjnnv|�������ztz|~��������xj|�̠j`lbL<:X|����zljnv~���������|vx������z�vjdp������jXV`jrxtv|�|vrv|������~ztx~���������||���������||��rb``bp����~��|p~���~|~xrt��ztx|�����xjjlv������~vdZ^ntvv|���������vt��vprljlnjlt~����z~�zh^h~���ztljv������jhz�zf\v������xFLhbj������~hRXz�����rRRjtr��������lPRhtxx�������z|�����xtplljp~������vjlnlfdlxxx��������~vz����������~�xh^`jrpnn~���������n^``bjttr����������vp���hV\x���fHRdt��������hZZ`TDN��ެf^���pLR|�����np|�����ldjdZXPHf�ξ���rnZ84X|����������t����RJX`bNLf���ʪztxT2^|�������Ғjx��lPLd~�������κtTtxF&(N�������zJJZX>@b�����������`J^hVFBRx��������vRJ8..D^~������ƒ���N"(DXZbbv��Ը�����f>8:Bb��l��¾��zppX,,J^lz����������zxnnhXTj�������ļ��XDNNJXn���vbTb���zf|�rB0HndZl���ή�vv���z|���vZR\z�����ƢrTVpfJB^~�������pLDRl�plx����|���������trz~pPFT����p��j0&<`����¼����~VBH`npv��zr���Դ�rp~h4&D`|���������`JLLPX^l�~�����Ҷ�|fF2.0:Jj�������ʠtv�zZ6(HVN\r�����ľ��X6.:N`hhj|��м�����rNJTVZhz���������`HJZjlbXZr���̲���|dN>Fd���ln�Ʈj���j<@P~fXP`p���ں�̚fB 4BDPh���ʪ����vF<VbVR^ft���������|f^Zdplv����������n@&8TPVp����Ғ���|N2<V`^TN\~�����ȴ�T8BTRN^|���Ȥ���pL>Pft���~v���������vR:2@JRb�����Ʋ��jTRVjtrb\ft��������x`PJRV`|��������xlnjhptlhhnxx~�������jRD@HXt�������~fZVZbnz���~���~�����ZVhr\JFTv�������xh\T^nxrdZh��������zffjj\HHh������Ĭ�ldjthPDNd~������������`RZbbZXXj���������hZhphfn������vz�ִ`Fr�t>(P����������ldvvh^j����h\f����z~��tLD`|�������~��~|~xtx|~zvlfhpz�~������j^bjlnt|�����rp|���������th���lr���pZXv��������~dZ^dflln|��rjt����lp���h^lz���������zzvlb\^frz|t��Ψ|nz|zpVPdrz|tx|�������rf`bprf^l���Ȣ����p^TXfz��|vz��������zfTBBTdl|�����РvrzlVJHb~~pv|��̾����xZPVdvzpr|��������rN:@Vbdp���������zlhnf\bv����������~phfdfjt~zv�����jbr�Ɯb^��~Z@Rx����|����z`v|j`\Rn���zr~���~z��rZJJVn�|x���ܶ�x|vfR4.Hhx~�����²���xL8DVTT`t��������|pbX`prrx�znp����tjv����zhnz|zx�������trzxnfp|||~�����������zh``fhhr~�����vhfx���������tb\`lv~����������xtxv|xvpv��xv������zvtpfdr��������|rnptzzzz|zxx|~~|�����rnlp|��~z�����vv~��~~���~|zx~�|zxtrv|���������xbPR^jtx~����xz��~pnr����xlp���������vbRNT`t��������t`VV^hv������������zvn^VPN`x���������zllrtnddr�����������xth\Z\bv����������ttpbVPVdt||�������vprtvxz�����|~��|z~��vlbbht~������������`JPbdTBFd����ľ��xvfPJTn���������|px�|n`blttpnx����|�����jTRdt~|rv����������l`ZVTZn��������zrphb`bffjv�����������lp|�thhr����vz����rhhjf^TP\p~���������tphdddp���������~����xrjlpvz~������~||xpjhp|~xtt|���||����|tz|tpnrx����������|ztpnllptxtnz������zrjdTNVh���������xfZ`t��������ztrtxz|xplp��������pfjrprrr~����x~���xz����p^^p��~z~�����zdXVXd~��������tffhp|��������~||���������~|zx~��zz|~|zz������vnprx|������zZFNdjhj|����������~rrxzxphhpx������ztv|tjffr~���������~|vpt~��xlhlz�������t���|t��~tnnxtf^ft������zxpb\XTfvrlt���������|f^fhptvz�������th^VZj|���������xpf`dr||ldjpv���������~|thdp��~xtx����nnr������z���xrpt��znjjv~��������xlb^bp��������znjhhn|����������zxxvzxtpllprrz���������vVJJLLJPXbz����ȼ��n^H<B^zz|�����~z���l\drpdX`v����������~l\TZfptx~������~z|xnbdfpv|�����������vh`^ZZbp~���������~ztj\TXdnvv��������vljpl\LFLdz���������pf`^``jrx������������t\^nz�~tt�����~vz����plnrvtt|��~~������������|vtvtrv��������|rt~��zvx���������rf\XX\blz�������������rjjjffjpvz~����������vj`V\lz|����������~vrlttf`fv���������rbd\VTZhz��������xnjjnpv��������zpjr���|vvvpnjhn|���������zh\TT\dlv����������������vbX^bfjpx~���������xvxz|zz~���vlnnrppv~���������������|�~xn`XZdnx~���������prxxz~tZZn��zv����|�xlnbZl|����������|XF:BV\dr����������|vvt|xf`nv�|~�����~�����vxvtvxvvtz���tlhrv|~������~|zvrv~�����~~vhVLTdtxx~����Ƭ���zfTPTbhjlz����|�����tf`f����������tlrvvz��tfjv���������xpjjhb`br���������p`VVfz�������|~�����zvxzzxz~�������~vv|���vr|������|tnjfjlrv|������������n`^dlttvz����~����������hTHN\hnv���������ztrtz~���~�~~z~���zv��~nbbjnrv~��������xj\TLNbv��������rntxxz��~�����|j^\fnt�������|tjht��������jhlbbXPXp~��������znjlhfpnx���x|��|z|�zt|��������vv|||������~zvrtz������������pd`bdbdlr|���������~���tf^`nxx|����������|vtttxvtt��������~tllv~xtx~������~|zzvrpx��������vb\frrnlz���������|tjhrvvt��������|xvvxrjfr~����������rf``fptvxz��������~tv���hjx||vpr����|xvtz|~|�������~|rlrzthj����|����rhpz|~������znfdhjlrrx��������z��vljnx�������zzz~�������~z|||zxz~���xtvx|�������~~��tf`ftxnb`v��ذ�z��~n^dnpx���xx��~|�������~|vttp`Vbv~~xzztrpt�����������p^ZXZ`ffht������������~z|�����vhddb^\`l|����������������vlhjnf\X`r���������|xtrtvz~���xh^^bhnrx����������~|~������|vnjlrvvz~����|z~��������xl^V\jrpnlt����xv����xllx�����z���|tvzrvvh^dnv���������t|~xt|�xlnv�������vvz���vdv����~�����zbNHP^r���������tfhz�������~���hNPbrrdRb�����������zz|phtz~~xff��|fbp��|~���tp~�������~|���nbjrtrjp�����v��ԶfDVx~�|b\n�����lf|���~~~z�~jfjt����z����hfhfhn|������������|trvtplr|����������vjd`\htx|~�������xx|~zvn\TZflp~��Ȭvp��xdX^z����zx������|rtjhVLV^bv����������xjTTfz��������tjdhfht��������zvjp������zh^V^r�|p|����~tx��lZbv��vlp����|z�zl`Zf���������~n`VV`jr~�xxzpnrtrpz�������|pjhp�������zrlflnhl~�����|����tbj||vrvxrtzvx�������tvzphlrv�����������rNNfvz|vpx~�����~���r``hbVVbt������������~tttppprx~���������zllppln~�������pdZV`d\Xdtz�����~���������|rp\NVf|��������|fpxlhd\bx�����rnvtfNNdrz����������rbflrnbjtvxz�����������fVn��fZr���|v����vth\z���bj���~j`hplh��������|lpnd^\`v�������rrvrnhnvxtpv������������phfnx��~ntz�|njhnxz�|zvtz���������zvtnbXXdr������Xl�ҔPJn��vVRz����������dPV\HJbr������֜v^`fXNLN^lvv����������xt~�����zxnnvnlvtp|���|rnlrz����������rbdjnnhl���������jP6,L��vNz�pLJ���~|����pTJ>L\f����������^D\~��np����pR\rjPZv��z~���������n`bVTf|�������zxxz��������~ttzzvv������lXVZ^`ht��������thht~�z|������~vpnpntz�������|rpt|�����~��~zzvptvxxz~��������~vx���px���|j^j|zndnzz��|xrrxtr������v���Z@Tp�zv~�����vn���tp����rt||~zhVZn���pz���������|z~�xpjp~~rjpz������������ztrlnrplhjpz�������������vpljhb`jx��������|jfr|���������tf`flnpt����|���~vv~�������~xtx~��|zz|~xrljnv����������|���rd^blhhpx|����vfd~���|�����z|�tZJP^`j|~���������nt�����thnpnnvvp~����vrndhx���������rr~�|vv|��rdp���������|pljjt|~�������zlddddn~xpz���������zvlbXLN\npz����zz���xz�����rh`Zbptv|����vf\Zj~rr��İ���vtjbh|������thtxdPX~��~l�����lt��~bdvzphhjnf^pvpz�������������p^RH>>JT`~����~���rjr|�������zphjv�������j\\`dn~�������xnfbdtzvz������~������~pd\VV^n�������zlfhlt~������x`RT\v��ʠ���~ZFHVr�������zphllnrv����zvrv�������v^RLPbz������z||vrpx|����tnzzz~����ƨr\\`\PLZ|�������xl\PRfz����|z|tb`�������zrdZVbv�������~xpp|��������zpffr|xtv���tnrtttx����������~x|xvxxxxz���������tplprt~�������~tlnnpv���~zxzxrrt|���������vjdbdhhl~�����~ztpnt��������n^XZh~���������vlntvx~����~vpppv�¼�lz��l\PVj||njjl��̘x|��t`XVbr|����´���jVJ>Bx��dv������t|~rlprnt�p`l~����������hh��`DPjnlnpx��������rld\bx���������jbfpz�~~������xbXV\^`r���v���v^RRn������xpttlhlx������xtt�����|���|tljlv|~���zvvtpnrt~����xtz��������|phZTZdv���������ldlv��������|n`NJPZflx��||~����������zlfbbjnnt|�������xvvz���������|nb^djjntrlt�������������xjfnx|rdft~���~�������tptx����~z���zhZXbp~��zrx���x~��������tbZh~��~z�������~zttz|vrv�������znn|��j`ft��vpv��������~�~vp~�|hp���vj`n���|rllv�����������lfddhr~��������pnt����������~rnjbbhrx|��~������������|trplptvplhjnz���������~tj^\l�����|phhd`bl�������xppt|�������zn`VPZfnz����������������~rlh`ZZ^bjz�����������|j^\dr�������xdN>>Pj��º����~bPVbn|����~~vptx���������r\R\jpnr|�������ztrpx��vpz��~|���vvvtx��������pbZbptt~�����zphb\h����������rjfdfp|�tln�����������vph`djpx|~�������|~�����|plljjjnx�������pd``fpt~�����~����nhr�vj`l��������||zzx�������zvh\Zd|�������|`VZbflv�������nXTl���x���~b\frndh����zn`j���rht�����th~����t|~dHBThlnv���ĺ�Zh|����tx���pVDLXn�����������xnd^fz��vljx���vhlv���zxz����������xvz~|tt|���znhjnz�������|tlbXPLVj|���������ztv|vtz��~xplp~��������xZRXbnrpx||~ztz���������`NJLRXj��������~l`b`\x���`b~����rz���xlbVP`ft�����������X6b���`NR~�|fhnz����z�����r����jLRp�~N8F`������������znlf^bz��zpl~���nn�����xvxz~����������xj`\\blx��������zt����xxxxrjbfpnfhv�����|�����rn|��xXBXt|ztv���������zv|����tbdv��pdl�����zxzzvvz�������~p~��rv��~rlhv��v�������|vln����x���zjj���h`rxzp`jvz|�����������pt�|^P^rx~xrrvx~���������Ȫ��h^PND<T^hx������������xjfrznrlbj����z����ptvvr|~������������ZL`vrhjdl����������vlfdx��rn�~tjb\h��xz������~|�����~z�~tf\Zh~�xrz���������~~���~xtrjddj��~v������vptpjz����~�����|rbdhjfhjx�������||l`^fr~�~z���~prx��pjv��zvvrjr~���������xddb\^dt���zp~������������\@:Pr����������vdZV^ntztrv|����v~����nfdbdhr���������v\RVZbr|~z�����z|�������xnhptppt~��������|zzxtppx~���~~~������zvvvvrrpx�������~~��znffnrvxvppv�����������vplfdp|�������~nhn�������~pjfhhjnv~��|vz�����������vfhnnld``l���������zx|�~b\p���|pn|�|rv������|����zr|~phhl|��xnt���znz��������zzxx|td`p�����������xtvtx~���zvtrtvx|~�����|xz~���|xx|���|zxttz��~||��������xz|~�~~|xprrtxz��������~xvtv|�����zvxztnjr|�������~vpx���~rx��zlfjx��~����~��~����|nrxxtx����xx~��|lj~��������xnr���pdjx��~xtt~��������zttprjht��������~vz~~~v|��������|xtrttxvzz|����~~������||||||z|~~�~����������~xvvvxzzx|������~xvrpnllnrvxz~�������xvld`dpz��������������~xrtx|~����~|~��|xx|��|ttvxz~�����zvtv|���~���������������zttx||zzz||���~��zvtvx~��������|xttvx|����������������|~|~|ztt|���|~�����z|~�~zxz|����~||~~�~xvz��|z|~���������|xtrt|����|~���vrrx|xxtppttx���������xhdp��xt������|~��th`dpz������zz|~xnlrz|zrv����~������z����~zzz|��������|tpppnnptz��������������vnljjjfhpv~���������~p\V`nxzz�������~|~zvnjrvz|��|z~���zrx���|txz|zz~���������|tlhnvz~����������zvrppnptx~~��~~zvvz������|���vjjpz~��zx~���������tvx�����~rx���rnt���|vz~�~�����~zxx~~�����|~�|||~����|�������~��~~zx|���~~~|xvvxvz||ztrpz�����~~���zxz���~xtrvxvvz������������zvtxz|~�����|xxxxvz������~||zxx|����~|~~���~zxz|||x|����|zxxxxz�����������~zzzzz|~~~~~~||z|~��������~zxxz|||~~||||~~|zxz�������~��vh`bnvz||������������vr|���|f`lzxl`dz�������~vlfhx����z~����phjv||vr~������|tpnhhr�����t|���pjr~��������|tnptz���������j`fnvvrtz�����������vnnz����z|��~vrx����~ztprvphnv~���������zz||~||~�����zvv|��������|zz|������~zxvvxx|~~zz|��������~zz~�������~xtrv|��������|zz~���zx|�����||zxrnnt|������|ztnnv��������~vlhlpvz~~���������vnpx�����xvz~zvzz�������~rlpz��ztpr|����zxvvvz~||������|rptzz|����~������|~�������~|xtnhlrx|~��������|���vnnv~��ztrttrtvz������������~~��|trv|~~xxz|~������~~~~�����~����zlhpz~ztprz��������~xtz��~nn|���xjl|�������~|vttprpjjr����������vjpz����|vxzvtllprx����������|pfdfjpvzzz|��������������vnlt|zxvt~������|tnpz|vz������|zzvppx���~�����~vvz���~�����~zvx||~���������|xvtpptz����~|xpr~���������h`dnpllnp~���������zlhp���vv����tlt���vtz|||���~||~|zzz~���zxxxz|~�������|z|xtx|�����~��~zxxzxvvxxx~������xvzzrlrz~����|�����������xvz��tjhjrxzz~�����|zzvvxz~||�|����������zz|~����~||zxxz|���~zx|~�~~�����|z|~~|xvz~�������|zvrppx~��������������������|vpnllprx~�����~z|�����~xxvplprvvx|~������������~���||zxjhpv~�������trprz~��������rllprrrt~�������~z|���������|tlhhjlr|������~zvrv��������|tjd`bjrz�����������������~phhfhhhnz����������||���~vnnpppppv|��������������zxvvz���|tpnrx|���������ztx�����vntvvfflpt|������x~������vx���pXVV`npt|���������zxz����vjjnvvprtz�����������~zxxvrtxzzzvrrtz~�����������~~������|trpnpprpnp|��������~vh^`hr~��zxxvrx������|~����|ljpxvnnz�����~rrvz�������zxx|�zplnv|���������~|z|~����~xrrtz����������~zttxz||~��������xxz~��zvtttrnrx~��������xvx||vpllrz��~||xvx|����������xnfdhnrx~��~�����~~�������~vnpv~���||���ztpnnprrv��������xjbXXhv��������rr|�����������vdZV\`dp~�������xppz�������|z|tphhlt~��������~zrvvx~�����|tttttxz~~�������~tpllnpxx~�����|xvz�����������znhdflrx~��������~|~����|xrprtzz|��~�������~~|��������������|xz���zxzz|���~|~������������~zrnpx|����������~~~|~~||zz~������|||||~~~||���������|xtpnlpv~��||z|������~|~����~|~��|zxxz|~����zz~�������~|zxvvxxz~������~���~|��������zrlfhlrvz��������������������~xpljlnx��������|zxxz|~|||xvv|�����~xx||xz~|zxxzz||~������|tt|zz|zrljtzxvzxz������������p^Z^dhlt~��|��������������vjhhd`bdhrz�����������������~xn`Z\^fjr|�����������������~pfddddfjr|��������������~~|xvtnhfhlrx~������������|z|~���~xtrpppptx���������������~|||zxvttttvx|��������������~|xtrrvz�����|zzzz|~��������������|ljnrnp|�||~������z|~����������vjfhjnlr~�������������������xttrldfnt|��������~~�����������vrljhlrtx��������zvvz�����~||zvplhhnv�����������zvvx|����~|xvrrrpnpx~����������~~~|z|||zvrprv~�����������|xz|~||�������~vrtz�����~||~|zxz||���|vvz~����zttz~�~|xrptz����������thbl|�����pv|�rdlpnv�����������vjlvz����zjrxrnhlr|��������~~zttrv������|rjfdfjt~�������|xtvz|�������zpjfddhr����������|vtx~���~|vrrnnrv|~����������|z|zxvxxvx��~z��zv���~�������|xz~~�����|������|ppx|�~|~����������~~xrlhflt~����������|zxz���~zxttx~��������������zvtppprz~��������~���|z|������zrprrrttx�������zxxz����������xnhfhlrz�����������zrtz����xlhffdblz���������vjjljnnrvx~�|z|������������vnlfbbfpz��������|||~��~�~����xpnptz~��������vpnllpv|��������xtrprv|~~��������������~~~��~xlhjnxxvz~��������������~rnpptvxxxz������������~zzzz|~����������|vrpnnllllp~��������znd`jllrx�����|z�������������rlf\^Zbpx~�������~|z|�~~|||~�xrjfhlv|���������xpljlpv|�������|xx��������ztld^^bhp|���������ztnhltz����xnnlhfp~���������~rljlnpv|�����xvvvx|���������zrpljnt~�����~xxvrptz~�������~vvvvxx|������vjjlprx��������~vrppvz~��������~xttv|~����������~������|tpnnlptxz~�������~|~���~|~~|xvtrnrvz~����������~~~~������~ztttttvz~�����������~||xttvvvxxvtrtz�����������|vttrtx||xxzzz�������