��������������~����~}~~~��~~~}}}}}}~~~||}}~~~~���}{{{|}}}||{zz{{||}}}~��������������������������}{{{{{{||{{|||}}||}}}|}}}}}}}}��~}}}~~~~��������������������~~~�����������������~~~}||{{zzz{{{|||||~������������������������������~~~~~~���������~~~}|}}}}|||||||}~}|{zzzzz||||}~~~~~~}|}~~~}||}~���������������������~~~}|zzyyyxyz|~�������������������~~}|||{zz{|~~�������������������~}~~~|{{zzyyzz{|}~~~~~}|zz{}~~~~������������������������������������~}{{zzz{{||||~~�~����~}|}||zyxxyyz{||||}}���������������������������������~~~}}||||zyxyyxxy{||}}}}||||~���������������~~~~~��������������������}|}}~�����~~|ywwwxz|{{zzz{|{zzzyz|~~�����������������������������������~~}{|~����~�}~}}}{zz|~�~|{zzy{|{|}|{{|||{{|}~~}}~���~~|||}~~}~��}~�����~~�����~~~~~���~}}}}|}~~}}}}}~}}}}}~}}~~~������������������������������~~}~~�~~}{|}~~|{|}}}~}{|}}~~~�������������������������������~~~~}}}}}~}|||}~}}}}|||||}~~~~~}|{{{|}}||}||{|}|||}}~~��������������������������������~~~~~~~}}}~~~~~�~~~~~}~~~||{{{|||}~~������������������~~~~}}~~~~~}}}}{{{}}|{{{|||}~�����������������������������~�}}|||~~|{zz{}~~}}}}}|}}}}}}~~~}}||}||}}|{{||}}~~~��������������~~}}}}}~}~~~~~~}~~~~~~�~}~}}~~~}}~~~}~����~~~~~}}}}}|}||||||}}}}|~~~~������������������~}}}}|}~~�������}~�����������~}�������������������������������������~~}~}{{||}}~}}|}||{z{|}~~~}||}}{{zz{|}~}}}}||}~��������������~}}}~~��������~~~~~~}}}~}}}|{{{|{{}~~~�~}~~�������~~~~�������������������������~~~}||||||}|{{{zzzz{~~��������������������������������������}~~~~~��}}|}}}~~~}~}}}~~~~~~~~}}}~}}}|}}|{{{}}~~}|}}}|~������������������������~~~~~~}}|{{{||||}||||||}~~~~}|{||}}}}||||}}|||||}|}~�������������������������������������������~}||{zz{{{{{}}|{{|�����������������������������~~}}~}}}}}}{z{}~~}}~~���������~~}{{{{{{|{{{{{|||}~~~~~~~~}}||~}|{}�������������~~~����~}}||{zz{{{||||{|}~~�����������������~}~~~~}~~~~��~}}}||}}���������������~~������}}|}|||}}}~���������������~~����������~~~}{{{|}��������������������������������~~}|z|}{{}~~~|zz{|}~}}}}|}}}|{z{|{{|{{~~�~����~~|||||zzz|}��������������������������~}~}~~~}}�~~~||{{z{{~~~zxwwz}~~}}~}}{yz{{}~~~~}||}}}|{|}~�������������������������������������}}|}|{z|||z{{}|}|||~���~~~~~~|}~~}}~~~~~~~}}}~~����������}|||||}~�����������������}}}~~~}~}}~��������~���~~~}|{{|}~~}}~~}|}~~~~}}~~~����������������~~}~~~~�~~~�����~}~������������������������������~~~~~~~~}|||}~~~~~}}}}|~~�~}~~}||��}~��~}|{{|}~~~~}}~~~~~~���������~�~~~~}}}}|}}}}}}||||}}}|}}|||}}~~}||}||}}||||}~������~��~��������������������~~~|}}}|{{{|}~~~~~~~}~��������������������������������}|||||||{{{|}~~~}|||~���~~~~}~}}}}|||{zz{|}}}}~}~}}~��������������������������~~��~}||||}|||||||{zz{|~~~~~����}}~~~~}||}~}}}}~�������������������������������}||}~~~|||}~}|}~�������������������������������������~}~���~||}}}~~~}}}}}}}}}}}}}|||}|{{zyyzzz{{{|||{|~~~������������������������~~�������~~}~}}||{||}}~��������}}}~}|||{{|~~~�����������������~~���������}|{}~~}}}}~~~~~��������������������������~~~~~}}}}}}|||}}}|{{|||}~��~������~}}|||||}||{|{{{}~~�������������~~~~}~~~~��������������������~}}|{{|}~}|}~~~~~||}}}}}}}~~~������~}|||{zz{||||~~~~~~~��~~}||}~~}}~}~�����~~����~�������������������������������~~~~~}}{{zz||{zzz{|||}}}}~~~||}~}||}~����~|{|}}~~}~~~��������������}|||}}|{{{|}~~}}}~������������~~~}}{yxyz|}}||||||||}~~~}||}����������������|{|}�������~}|~~~~}{yxwxz||{{zz|}}|||}�����������������������������~~~}~~~~~}}~~~����}yxxyz}}}|ywwz|~}{zyyzzyyz{{zwuvxy{{{z|}~��������������������~}}}}��������������~~~}|{{|~}|||||{{|}|{{||{{{{|}}||}}}}~����������������������������~�������~~~��~�~}}~�������������������������������������~}|{{|{{zz{}}|{{|}~~~~~~}|{{{{{{{|{zzzz{|||||}~~�����������������������������������������~}}}|{||{zz{{|||{{{{|||}~~~��������������������������~}~~}}||{{{{|}}}}}|}}||}||}}}}~~~}~~������������������������������������~}|}}}~~~}|{|||{{|||||||{{||{{|}{{{|{{zzz{{{{{{{{|~~��������������������������������������~|||||}|||{zzzyyz{{{|}}}}}}}}}~~~~~~~}~~~�����������������������������������������~~~}|{|}}~~~}|{|~�}|}~����������������������������������������~~}||}}||||}}|{zzzzzz{||{{|}|||}��~���������������~�������������������~}}~~|{{|||{|{{{|}~~~~~~~~~~~~~~}|||||||||||}~��������������������������~~~}{{|{{||{{{z{}|{||~~}}~~~~������������������������������������~~}||}}}}||}}~~~~~}~~~~~~~~~~~}||||zz{|}~~|{z{|}}}~~~~������������������������������~~}}~~~}||{{zzz{{{|}~~~~}}}}~~}}~~}~~~~��~~~~~~~~~~~~~����~~~~~~~~~}}~���}||~�����������������������������������~}}}}}~~~~|{zyyz{{{||}~~}}~~~}}||}|||z{|||{|}|{{{z{|}}~~}��~~����������������������������~~~~~}~}}|||{{{{{{{{{{{{{{{}}}}��������~~~}}~}}}}~~}~��������~~}||||||{|}~}}}���������������������}|{{{{|}~~}��������������������������������������������������}{zxxyzyyz||yvttuwzzxxyz|���~~���~}~~}}}}|~���������������������������������������������~~~�~~~}{yz{zz{|}|zxwwxyz{{{{{{}~����������������~}|{|}|}~}||}}~����}}~~����~~�������������������������������~}~~}|{|||||{|}~��}}}}~~~~~}|||{z{|}|{|||}~}{{{{|}}{zyz|~~}}�������������������������������~~~~}}}}}}|||}}���������~}}}||||||}}~~~~~����������������������������~~}}��~~~�~}~�����������������������������������������~~}}}{{z{z{|}}}}}}}}~~~~~~}}|||{z{{|zyy{|||{zz{{}}~�����������~~��~~~~�����������}|{{{{{{{{{{yxxyz{}~}}}~~~�����~}}~}|}~~~~~������������������~~~~~~~~~~~~~~}|||||||||}}�����������������������������������������~}|}}}||}~~~}|{|}}||}}~}}~~~~}||}}~~|{{|}}}}}|zz{|~��~}~������������������������������~~}}}||||||||||{{||||||}|}}||}||{{{|}}}}~~~�����������������~�����������������~~~}|{{{}~~}~}}}}~~����������������������������������~~~~}|}}}}}~}}|{{|}~~��~~~}|{{||}|{zz{{|~~~|{{{{{}~~~~~~~~���������������������~~~~~~}}}~~~~~~~}}~������������~~}~~}}}}~}}~~}~~~~}}}}~������~~~~~~}|||||||}}}|}}}}~����������������������������������������������~}||||}~~}}{zzz{|}~~}}|}}}}}}}|||{zzz{|||{{{{{|}~~~~}~~���������������������������������������~}||{{|||{||{z{{{{|~~~}||||}~~~~}}|{z{z{{zy{}�������~}~}}|{|~�������������������������}}������������������������������������}|{|||{|{{|}}}||||}~~~}||{{zyyzzz{zzzz{{|{z{|~��������������������~~}����������������������~}||{{yyz{{{|||{{{|}�~|~������|zyyz{~~}}~��}|}�������������������~|{zz{{|���~||}~�������~~��������~�������������������������~~||}~}||}~~|{{|}|zzyzz|~~}}|{zyyz|}}}~~}||}~~~~}|{{{zz{|}}|||}~~��������������������������~}}|{|}~~~}~}|{{z{{||~~}}}|}~~}||}|{{{|{|}~~~~�������������������}|}~�}~������������������~}}|}}~�����������������������������������~~~~~~~}}}}}}}~~~}|}~}|||||{{{{zzz{{}}~�������������������������������������~~}|{|}~}|}}|{{{||}~~}������������~}||}}}}}}}}}}}}~����������~~�~~~~}}~~~~������~~���������������������������~~~}{zz{{}}}}||}}}~~~~~~~~~}||}~}||||{||{z{}}~~}}}}~~~~~�������������~~����~��~}|}}}}}|||||}|{|}~~~~�����������~���~~}}}}}|~����~~����������~}~~~~~}}|||}}}}}~~��~~~~~������������������������������������������~}|||}}~~~}}}}|||}||||{{{||{{{{{|||||}~}}|}~~������~��������������������~~}}~~~~}|{{|}}}}|||||}}~~}|||}}~~~}||}~~~~~~~���������������������~~~~~~~}}~~}|}~�������������������������������������������������~�~}}~~~~~}|{{||{{||}|}|}~�~}}}}|{|{{zz{|{{{}}~~}}~����������������������~~}}}~~���~~~~~}~}}}~~~~~}~~~~~~~~~~~}~~~}}}|}}}~�������������������������������~~~|{}}}}~|}~~~~~���������������������������������~}||{{zzzzz{{zzz|}~~}|{{zxxxz{{{}~~}}}||}|||{zz|}~~}~��������������������������������������������~}}||}}}}}|}}}}~~~~}~}}}}|||{{{|{{yyyyz{{|}~��������������������������|{zz{}~���~~~~}~}}||||~~~~����~��������������������������������~|||{{|zxxxy||{z{{||{{|}|}}}|}|}~~}}{zyyy{|||{|}}|{{|}��~~�������������������������������������}zy|���~{z{{z{}}||{zzyxwwwxxxvvvvvvvyzyyzz|}~~}���������������������������������������~~~�����~~������������������������~~~���~��������������~~~~}~}}}|{{|}}|{{{|||||{{{{|}}|{|||~����������������������~~~}}~�~~~~~~~~|||}|||}}~}~}~~��~~~~~}}|||}~}|{{|}|}}��������~�����������������������}}}}~�~}~���~}����������������������������������~}}|{{{zyxyzzzz{{{{|}}}}~������~||}~}|{{{zyyz{{{{|~}}}~��������������������~~��~~}}}}~~}|{zzzzz{{zzz{{z{z{|}}}}}}~~}}~�������������������������~~}~~~~~~�}~�����������������������������~~~~~~~~~~~��~����������~||||}|{zyyyxxxz{zzzzz{}}~~~��������������������������������~~~~}}}}}}}|||}~~}}|||}}~}}~~~~~~~}}}}|||{{||||}}~�������������������������~~~�������}~~��}~~~���������������������������������������~~}}}}}|{z{{|{{{|}~}}|||}���~}}}}}{{{zyy{{{{{{}~~����������������������������������������~}||{||}}|{{{{z{{{{{|}}~~}}~~}}}~~~~}}}~���������������������~}}~~~�������~~}|||}|||}{{}~�~~������������������������������������~}}~~~~}}~~�������~~}zxyyxwwvvwz||||{{|}}|}|||~��~�����������������������������������}{{z{{{{zyxxz{{z{zzyz|~���������}}|{zyxxyzz{yyz|||}~���������������������������~|{|~~~~}}~���~}}|{{}����������������������������������|{{|}}}|{{{|}~~~����~~}}~~|}}}|{z{zz{{zz|||}~}|{|~}{{~~}����������������������~~~~~~}||}}|}~~�������}{zzzzzywvxy{||{zz|||zyzz{|~��~������������������������������������������~~~~|}|{zzzz{|~��������������������~}~��}|{{}}}|{z|||||~}{yy{}~}}|}||}~}~��~|||}}~~}||}|{zyxyyzzz{|}~���������������������������������������������~|{{z|{{{{{|||{{{{||}}~~~~~~}}~~~~~}}}}}}~�~~�����������������������~~���~~}||}}}}}|}}}~��~~���������������������������~~}|{|}}}~}|||||}~�~}}~~������}{|}}||||}}{zz{{{{{}�������������������������������~~~~~|{{zzz{{{|||{{{}~~~~~~~~~~~}|||}~~����������������������~}|||||}|{{|}~}}|}}~~�}||{zyz{}}~���~~~������������������������~~~}~����~~~~~~~~}}}}}}}}}~}|{zzz{{zxxyzzz{|{|{{|~~~��������������������������������~~}~}}||{{||||||}}}}~~~~~~�����~~~~~}}}}}}}}~~}}|}}~~���������������~}}~~}}|~~~}~~~�~��~~��������������������������������~����~~}||}|{{||{|}~~~}|||}~~~������~}}|||}}}~~||}}}}~~�������������������������������~~}||||}}}}}||{{{|}}}}|||}}}}}||||}~~~����~~}}}~~~�����������������~}}}}}}}~~~}}~��~~}||||}~|}������������������������������������~}|{{}}~~~���������~||}|{{{zzzyxwwy{{zzzyyz{}~~~~����~~������������������������������~~~~~}}}}}}}||{zzz{||}}�������~~}||||}}||||~~���������������~~����������~~~}}~~����������������������������������������~}|{|}|||{{z{{}}~�����~��~~~~~}}}||||||{yxxyy{|}}~~~�������~~������������������~~~~~~}}}~~}}}|{{zzyxy{|{{{|}}~~����~~~~~~~�~~~���������������~~}|zz{}~~~~~~�~~~�������}}�����������������������������������~}}~��}zxy{}}|}~~~}|||}}}||}}{{{{|||{{{{{{|}}}}~}}}|~~�~~�������������������������������������~|zxxyyyyxwvvvuvwyyyz{|{yz{{|{|}~~~}}~��~}}}}}}}}}~}|}~~~~���������~~~�~�~}}~~����~}��������������������������������������������~~}}}|}}|{zzzzzy{{{{||}}}~~~~~~}||||||||}||{||~������������������������������~}|z{{zz{{{{zyzz||||||}}|||||}}}}}}}}~~~~~~������������������~~~~~}~������������������~~}||}}||}~��~}}���~����������������������������������}|}}|{{{{{{|}|{zz{|}~}|{z{{{z{{|{{{{zzzyyz{{|{{|}~����������������������������~~���}|||{{{|||||}|{{||}||||||||}}|{{|}}~~~~~~~~~}}~~�������������������������~~|||}~~}|{{|}~���������������������������������������������~}|}}}}}|||{{zzzzz{{|{}}|{{zz{{{|||||||}}}}~��}}���������������������������~~}|{||}~~~~~~~~~~}}}}|{{|||{|{{||}~~}}~~�����~}|}}~}~~����������������~~}~~~}||||}}|}}��}|~~~��~}~�����������������������������������~}}}~~}}|}||{{{{|}~���~~~~~}|{{|{zxwvwxyyy{||{{|}~~~�������������������������������������~~}||}}}||{zyyyzzz{|||}}}~�������������~}||||{||}}~}~~~~}}~~~~~~~}}~~}}~~~}}}~��������������������������~�����������������������������~}|}}||||{{||}||||{{{{{{}}}}}|||}}}|{{||{|}}||}}}}~~�����������������������~�������~}|}~~}||||}||||||}}}~~}}|{zz{|}}}|||}}}~~~~}}~���~}}~������������������������}||}}|}}}~}}}~}||}}��������������������������~~~}}~�~}}~~~~~~~~~~�����~|||}||{||||||}|{z{||}~�~~��������������~~~~~~~��������������}||{z{}~~}{{{}}|{|~�����������~~~~}|}}|{zzzz{|}�������������������������~~|{||{zzyz}}|}~~}������~{{|{{|~�~||||}~�����������������������~}}|zxy{||}}|||{|}|{|~�~~~}|~~~|{|{{||{{|||{z{}}}������������������������������������������}||||}|{{{{||||{{|}}}}}~�~~~}|}}}}}~~~}}}~~~~~~}~��������������������~}}||{{|}~~����������������������������������������~~~~~~~~���~}}|}~~~~~~~}||{|{z{{{zyyz{{{||{|}~~������������������������������������������~}|||||{{{{|||||||{{{{|}}|{{{|}}~~}}}|||}}~~~}}~~~}}}~~~}~~�����������~~~���~~~~||||}~�~��~}~���������������������������������������~}}}~~}|{{|}}|||}}~~}~~~}|{{{{zzz||{z{{{zyz{|}~~~~��������������������������~~}}~�����~}~~~}|||{{z{{{||}}~~~~~~~~~~~~~~}~~����~~~���������������������������~~~~|{zzz{|{{|~�����������������������������������������������������}|{{{{{zzzz{{{zzz{{{zzyyz{||}}}}�����������������������������~�����~}}||||{{{|}}|||}}}|{|}}}~~~}}|}}~~~~~}|||||}~~��������������~~~����~~��������������������������~~�������������������������~~}|zzz||{{z{{{||}}|}|||~~~}|{zzz{|{{|}}}}|||}~��������������������������~~~~~����������~}}||{||||~~~}|{||}}}}}~~~}}}|||}}}}~}~~~}~~~~����������������������~~}}}}}}|}�~~~~}}}~~��~������������������������������~~~}|{|}}}}~}}}~~~��������~~~~~~~|zyyyxxyzzz||}}~~}}~������~}|~�������������������~~~}}~~~~~~~~~~~}}}}}|{{{||||}���������������~~}|||||}}}}~~~~~~~~�����~~~�����������������������������~||{|~��~~}����������������������~~}|}}}�~~|zz|}~������������������~}}~�}{~���~}|}~������~~~�����}|||{{{{zzzzzzyxz{||zyyyyz{|}}}~~~|||~}}|{{||}}}}~~~~~~~}~~�������������~~~~~~}}}}~������������������~~||{{||{|{{~~~���������������������������������������~~~~~~~~~~}||||~~~}|{{{|{{z{{||||}||}����������������������~�����������~~}}}|}~~}~~~~~}}~~����~}}~~}|}~~~~~~~}}}���~~�����������������}}~~~~~~~}~~~}}|}}}~��~~�����������������������������������~}}|||||}}}}}~~~~~|{{{{||||{zz{{{{z{{zz{||}}|||}}~~~~~~~~���������������~}~~}~~~~~~~~~~~�����~}}~~~~}|}}}|}~~~~}|||||}}||{{{}~~}}~�����������������������~}||}|||}}|}}}�����������������������������������~~}}~~~~~~}}|}||||{{{{zzzzzzzz||}|}||{||||}}}~~}{{{|~~}}���������������������������~~~~~~~~~~~}||}}}~~~~~~}}}}}}}}|{|||{{||||||{z{{|||}~~~}}~���������������~~}}~������������������������������������������~~~}||||}}|{|}~~������~~����~}}}}}}}|}}}|{{|{{|}~���������������������~~~�~~���~}}}~~~||{{{{|}~~���~~}||||||{zz{zzz{{{{|}}~~~~~~~���������������������������~}||~~}~�������������������������������~~~~}}|{zz{{||{{{{|}��~}}}~~~~~}}~~~~~~~~��������}|}~~~����������}}~���������}||{{zzz{||{{z{{|}}|||}~���������~~~|||||||||||||~~~~�~�������������}|}||}}|{|}~~~~~������������������������������������������~~}~}~��}|||||||}}~�����~}}~~~}|}}~}~}~�~}}~~~~~��������������������~{{}}|||~|{zzyzz{zyyy{|}}||||~~}z{|}}~}~��~~}}}~�����������������������~��������������������~|{|~�����~|||}~}{}~}{{|}}|zz{{����~�����������������~~~}}||{z{|~~}}||}}|}}}}}}~~~}~}|{{{zz{{{{{|~���~~~��������������������������������������~~}}~}}}||{{||{{|{zzzz{{}}}~~~~~~~~}~}||~}||{{|}}~����������������������������~}}|}~~~~~||}~|||{|~��~~�������������������������������~}~~~~~~~~~~~}||}|||||||{{{{|||{{||{z|~~~}}~�������������������������������~~~~~~~~~~~~~~~}}{{|}}}||{{{{{{z{{{{{yzz{|}|||}|}}~~~~��������������������������������~~~~~~}}}{zz{{||~~~�~~������������������������~~��������~�~~~}||||{{z{{{zz{{{{{||{{{}}~|||{{{||}~�������������������������������������������~~~~~~~~}|{{{{{{{|||{zzzzzzz{{}}}}}}}}}|||}~������������������������������������~|}}}~~�������������������������������������~~~~}}}~}~~~�����~}}~}}}|{zyyxxxyz{||{|~~��������������������������~~~��~}{z{|||}~~~~~�����~~��~}}~}}}}}}||{zz|}}}}||||||}~~~���~�����������������������������~}}||~~~~~~�����������������������������~|}}~}}{{zzyyz|}}}}}|}~~}~~~~~~~~}}}}||{{|}|||}~~~������������������~�����������������~}|||{zzyyy{{|{{{|||}~}}~~������������������~~~�~~}|}|{|}}~~}||~~}~~~}||{|{|}~�������}~~}~~}~~�����������~}}~~��������������������������}}}}|{zz{{{{yyz{{||}}}~}|{|{zz{z{{||||}~~}}|{z{}�������������������������~~~~~~~}|{zz{{{z{zzzz{{||}}~���������}~}||||}}~~�}~~~~~~�������������������������������|yxxxxy{z{|}|{yxxww{|{}�������������������������������~}|~�~}~}}|}~}|{{zzzz{}~}}|}}~~~}}~~|}���}|{{z|��~~|{z{{}}~~}}|||}}~~}|}~������~~~}~}}~~~~~||}~~~~���~~~~~~|}~}~�~~}}||~��������������~�~~~}~~~~}}}}|}~~~~~}~����������������������������������������������~}|}}~}||~~~~}}}~~~~~~|||||}{zyz{||}|}{||}}~~��������������������������~~~}~~~~~}}}|}}}~~}}~}}}~~~~}}~~~}~~~����~~~~������~|}|}}}|}}}|}}}~��������~~~~~~}}}}|~~~���������������������������~}~~�����������~~~~}~}}|zzz{yyzzyyy{zzyyyyyyzz{{|}~}}}~}}}���������������������������������������~}|||}||||{z{z{z{|}}~~~~�����~~}{{{{zzz{{{zyzz{|~������������~���~~����������������~}}}�����������~�������������������������~}{zyzz{{||||||||}}||{|{||~~}|{|}}|||||zzz{{}|~~����������������������~~�����~���������}}}~~~}}|||{z{|}|{zzzzz|}~~}}}~}}}~~~~~}}}}}||~~~~�����������������������~~}}}}}}}}|}}}}||}~~~�����������������������������������~~��������~}~~~}}}||{|{|{zz{{|}}~~}}||}}~}}}|{{{|||}}}~~~���������������������������~~}}||||{{{|||{|}}~~~}}||{||}}~}~}|}}|{|||{||~~~}}~~}~~~~~~~��������~�������������������~}}}}}}����~~}}|}~��������������������������~~~~~}||~����~~}}|{zy{||||||}~~~}~~~}|||}~~~}}~}}}~~���������������~}~�����������~~~~~}~~}~~~~~�~~}}}}~~}||||{||}~~~�~}}|||||}~}~}~~~}}}~��������������~~}}||}}}~}~}|~}||}}~~~������������������������������������~}}}}~���~~~}������~}|zyxxwxvxyyxyxxx{~�����������������}��~~~������������}}}~~~}|}~}|}}}}~~������������������������~}}}||{{z{{{{|{}||{}~�����������}|}~�}}~~}~~}~~}{|||zzyz{|{{{{{}~}}��~�����������������������������~~}~~~�~~}~}}{{{{z{{|}}|z{|||}||{|||{{{}}~~}}~~~�����������������������������������~~~}}~~~}|{{||~����~~~~~~~~~~~||{||||}}}||}~����������������������~~~}}}|}|||}}}}~}}}}|{{~���������������������������������~~�~~~~~�~~~|||}||||zyyzzyyyyyxxyz{{}~~~~}}~���������������������������������������~|{zzzzzz{|zzz{{||~~~}}}}~}}|}}~~}|||}|||||||||||}~~~��������������������~~~}}}}|{z{{|{z{|}~~~~~~��~���~~~���������������������������~~}||~}|{{|}}~~}}}~}}~���~}}}}||{{zyxzzz{z{}|{|}~��������������������������~~~~~~~}~}{{|||}}}|||||{{zz{||}}~~}}}}}~~���~~||{z{|}~~}~�~~������������������������������}}}}}~~}~~~}�����������������������������~~~~~}}~~}}|}|||}~~~~}|||}~~~}|{{{{||||}~~~}~~~~~����������������������������~~~~~~}}}}~~}}}~~~~~~}~���~~~~}|||||{zyyyyyxxxxyz{{|}}}~�������������������������������~~���}||~}|{|~~}~~}}��������������������������~~~��~}}~~~����������������~}|zz{zyyyz{{zyyzzzzz|}||~~~�������������������������~}~����~~~~����~}||}~~}}}}}}~����~~~~~~}|{{z{{|}~��~||||~������~~������������������~~~}{z{zyxxyzxwxz|}��~�����������������������������������������~}||}~~}|{zyzyz{{}}}}}}{{zyxyxxyz{{{{{{{||{{|}~��������������������������������������������������~~}|||zzxxvwxyy{|}}}|{{{{{||}~~}}~���������������������������}zxwwy{{|||{|||{|}���������������������������������~���}{z{}~~~~~~��~~~}~}||}}~}~�����~}||{{|}~~~|zxxy{|~}||||~~||~����������������������~}}}|{{}}~~}||}}|}}}~~~~�~~~~~~}}}|{zzyzz{||}}}}{z{|~����~~~����������������~~����~~}}}}|}}~}���~�������������������������������~|||~~~~~}}|{|}}}}}|~~}}||||}}}|{|||||{{|}}}}~~}~���������������������������������~~~}}|||||||||}}~~~����������~~~~}}~}||}||}}}|}~~~����������~~|||}}~~~���������������������������������~}}��������}|{zyyz{|}}{{{zxyz}}|{{{{{|}~~}}{{{|{|{{{||~}|}}}}~~}}�������������������������������~~~~|{{|{{{|}|{{|||}~~~~~}}~~~~~~~~}|||}}~~~~}||}|}}~~~~~}~}~��������������������������~~~}}||||}}|{}}~}}~��������������������������������~~}}}{|}}|{{{{|||{|{{|||~�~~~~~~}}}}}~}~~~}}}}}}~~���������������������������������}}}~~~}}|}||||{|||{{|}}}}}}}}}}}}}}|||~~~|{{{||}}}~~~~}~~���������������������~~���~}}}}}}~~~~~����������������������������������~}{|}~~~~}{{|}}{||}~~~}|}~~}}||}}~~~~}|{zyyyyyyyyz{||}~����������������������~}}~}{||}|}}}}}|||}}~~}}|||}|}}~���������~~|}|{z{{||~~~~~�������������������������������}|{{{|{{{zz{}}}}~||}~~�������������������������������������}}}~~~}}}~~~~~~}}}}}}||{|{||||{{{z{|}}}}}}||||||}~���������������������~||}~~}}|}~�~}}}|}~~~~~~}}|||}~~~~~}|{zyz{||~�������~�������������~}~~������������~~~}}}}}}|||||}}}}|}}}}~�����������������������������������������~�~}||{{zyyyxxz|~}||}}}}}~�}|{ywvvwxz||~~~~}}}�������������������������������������}}}~�������~~}|{zzzzzz{|||}~}|||}}|{|}���~|yxvx{~����������������~~����~~}{{}}��~}}||}~~}||{{|}���~}�����������������������������~}}}}||z{{{|}~~~~~}~}~}}}}}|{{zzzzzy{}~}~~~~~~����~}}}~~����������������������~�����~}~~~~������~~~~~~~}}}}~|{{{{||||||}}}~~~}}~~�������~�������������������~~~~~}||}}~~�����������������������������~~����������~}{{|}}~}|{zz{|{{{||||||{{{{{{{}}}|}||||}~����������������������~~����������~~~~}}}|||||}}~}~~~�������~~~~}}}}}~}|{||||{{{||{|||{z{|}}~~����������������~~�~~}|}����������������������������������������~}}|{z{{{zzzzzzz{|}}~��~}~~~~~}|||}}}{{{|||}~�������������������������������������~~}}}}}||}~}}}}}}||}~~}}}~~~~�}|{|}}}||||||||}}}~~~�����������������~~��~���~}~~~~~~~}}~���~~�����������������������������������~~}~~~~}{{{|}|||}~~~~~~~~~}~}{{{z{||z{zzz{|~~~������������������~�������������