���Mʪ6������:�7�{��[����fq���D��s�.����a�9�_#�����ة5g�S�3c�p�Ȟ��^��s�cM��R�q�H��mJ��ķ�8r�ω�4!�i
�]����0%�1�i��݊�l���k�n�F��vS�_S���f%Xkæ]�ݎ3G1Y���e�uyu�B�������5���?O���K��:1���).>��DǿT�b�(t�[�X} _;<�ys8��8�	������~';�D2�Ұ��2���aus���R�Q�T ������tTZ����!R �_�%�~�#�����sZ�>^#'B�G����|�����?�3��g�'Y����?6*����A���B���*�������z /
v��T2��k�p��O��g��A�˝y��N������y�m0�g,��p��/Ć���"���H�I�lբ�a���	�y��&pD�a�����u��pw�}�rYhz'�}S�	q���ZC�V�*ژq~����(�"�9~�Q�Id'2����g)� 8:��n)�� j0Zh���`Z���������@����e�R�Ȯ��Wq���Z�>d��A�B��#����2=��V2O�*H���.�Of��o(�L�w*j�q�~k�1Q_)� �=�#3_�v�z{�wA���K]���wT[4�
 �~`h芬���R⪢D��{N�7	�f�c��דnh>Z����rJ�A+�wva�)T$����bExC�b=^�D��O-��V~?pс ��i��lK�@ÀccCF��f��)��z�~g��s���W
���G3f��Ѽxa��ʃ�+�P+Ѹb�KƥN,y:V1}��,qI}�e@R}�`-�r��e/qĝr��b�����'��K�Nb@ �B�+�f���F����f3;#_�VV�����IvE��v�ǜ<�<<�V�����hX���;�����(Q*�6r8�>,5���x��XZ�R�k�D1�Ť�J`���5����6m���Y�_�s���9u����B��$����0dZ�b�):��<�0fޅC?����k%��� Hv}��k�9��!�Ņ��b9o�cmU,g��eS���;��HD5,�ɹ��vj���������l�x?��k;+�"Mǻ��I =˿6:�5>˶�����]\U�v��iFz��%w�,��V�y[��*�����	��߆���]�9�Y��5��cU)g6o�3�71�|��skv���6�������:�� �%'�������?��i�NQ