�Dɔ5�߯p�R�M��zA����U�b�!���@�ӯ����f%��e�;)C�53V�[�܌��C�4[<�a�kL=�s��d$s�I��C8��*�~��9����9��O���k�	v�$c81J������{lt�u��SM����3yg�d,W�҉����v0!���Z�"�N?d�V(�f��Xv�^kf���J�tB5H�%���+69C4_8���V������:NCs���7u�q��+8<�	�B��~���Q�X}���������W��b�漭c�t��Ah���F��60��(_N��ݾd�x#�����Z��c�꥔���$ys����确:��p��̋�Y�6�؋��ȇFIc��[y 4�6ն�c`��珈BRaj��Oa��1����Q��H��>K����1����%��)��'��i0��a|(Ƭz姚�Pz��'&�I��?\��W��*DJ��AZOrV��L(��3W�34��V����eNq�[~��y���2��L��d>#�ѬP7�83y�dgY�e��%t�$��Z��IJ@.�/j��_ ����>ǅ����Z$���p8*ʡ��)�����O�*�bh��g�����k�X�,��#�$D�����KU���^�f��hH8�g�� f!h�]�Ĕ%�1�uf[�,0���E5�_�0�����n��9Ũ���w�%���j�����^4Z�?�3���`9C�1�ۛ�7"7/���^>�v�L7�p�IE�7���M �	|N�ϓ<��[������zдt�cny#�d���\����S �����#��@�����ǐg,�F%Ber�,!.ڝoM���P?Of�Ba�������L�B?��@@r���S��I]&�b��:�	P�B�dW�P�����x�y�$�͆�����w45 ����)�&n�3�F-������# ݯ�s ����ّgk��A��{��:����ň��cd�v&���bCz�&܊�Q�l��V9K�׆k��ߘ}7����H��mec�dX�En��t��$�i��P��P�嘎I�^�j{f�QD�a#�ɑ�h�kW$�qw�sX��ߪi@'�&���3��:�����#ǅ��OZ��aNa�ڻ����m��|�k�Su�QD.z+ZY��<��f�z"ueG}:r����P�T����F��T�ｻP�4�"���1��L	�G�c��Kò�! )U���{3{���(�<�ȡ\6X���#-͢�P�3���|U��qY*���m��B�M|>�$J8��8����k�2
��L�݀gq��� �vL�T�N׆��1�OEr�ĉ�΢��������tB|�L\/��-%}]���`��Lg�^�iMJxĨ�lf��8�BbB`9�/��/�f�+$���zwخ(�3��'?�3ɔe2BU�)v� mx����&�"!lL�:,?�:�y�~�{�M(`v�7���K�b�&E��[���\Ld`�Ҍ����?q�m��A$+�y+�#j�t����5�N��Q^Г�I[dB��c��B��L��i|1�IcH��l:�]���8�&/c��ڨc��X����̟e��<T������>��dcON�d���eפ�xQi�͹���嶐����]��v��}���.�$p���v�Q#%��)�r�l<����	����́8W@� �/�8�dS�\���5j���h-<r�
�����C��#�碛i���J����'0iN'W�����&��Ļ�+p���I�a�%�=X�6k�<1Ʀ-$���;9��$��t�pMk<�_�L���BPy�Qp|��d^�toU:�rؼېb�Z�AC :��B8Ʈ����E����5�!�O�by%1�](�2:��yh����-�?eprY��ʂ_<r�i�խV����lCG3v�=��&!�(���<W��u=f*^�Mh

zz����>#3�2�Y��RޱT�k��"RG�f�i@�F�آH�p��u��4`�m;|���7�N}���L�!���F�_�#�����ܑa��qF��s�������$2_G�7��IF�=+񔋝�&Pz��p��)1,�]Et3U�7>�͹_^�2\-%��-Yޒ�-u��ˑDU�bR���J���;�,[M�?��4�v&����f��kꩽ�ǟ�����g��65�'r��`+�n��|��u<ͨ��gP�P	��t���E<�HG,��:�a���%J�6K=cb(y1��֡
�؟�Z�����	�ԔcX>�[s����я�S��@a�oѓ�Z1a$�:�e�s���z�cx=����gO����҂�c�mI�y�bO?�d0��ɺB��j�@�O:�ߚ�-@S���QG����=�ac�,��:��a\��z�s-f8�Y2B����	�@:�r"���d�ni��u�QJ[� �Bm<���+��/A��Y�7���0�Dl\Mv�m�* �7�S(�[���x���Դ� 8�������R�B!;����l����Mt�ZL`�VA�Z ��n�7���S��A��@ "�Zz���u%A�h�2\S�L��� z������S�)l ��I��原i��o�\5����:��.˿'ϋ�������$'�44[X� '�v֠#��y����ޤñ�>B���Ş�
T7�t+<�cð��[�d�����u5J���N���p)h���T��y��dl8�z��D8ٝ�I�Ou�~�M��E�y7�G�=~X��y�F}0��>B�&��)B8h�}5v��>O����H�X�D�����g�a�/thR�{^bC��H&������v�'�����Ћ5:�@'&6�m�T#LgF�a+֬�����5����l<���c�(�������K�~���e[�������C�;p��4!U��R��п7�3
��L�h�a�m��gE�V�����O�]Y�N-!(l�a��!Y,�Ş�#Nx�k��d��r�rb�)
;�M� �#������'���?�m����K�dwT*�
�pu֟��������f���� �w�3��1[�ch��nO��KLM�˛_1�E���ؙ$�8�@հ\	F�C:E+�~���N�<�Q2D'L�Z�K�b�k9�O��zivUe��6I)�:�K�9�rR袚][��V���4F��c��.?"�ۑʤ~���a��,�S��L�����������,��l)�T�O�(3�Z=����cvSf�Yc&2��Y�}�O����z�rybv���p���\�.p[흹��i9-2����S
S����)�,�F:OiÍDL�!��t��|lr���^XJ���K��fe5�<6q�s$yͤ�]����b&?c��|��9ſN<������(�ω�N]n��|@���X �R��kxE1���v�=/6�L�߇i�6'�N�0!�`�Õ�j��4�R'y����]<�=־��o��ץ���Z	t%c�7z��ʝ,	�m�Ȍ��r�F�(	�)��(-�2^�h�ɣ�F�[Ʌ���B�,29�3�I�)���^ӍȾᐡ��fx_J�b�{�m�/_��&�+U��˷|4��Y�("%�G��kl��}��D4���	ns�9)�/�+m+�&������qE]c����v g�
����,��e��Ϟ�M���x���lCj/���T�Q2�ہ�R})�ܽ���Q6�2�Դ�V\��ǆ�	'�����ܡfw�=K��;G(���z�*h���ޭ���q� -[�K�a4n�]>��z�;h�g w�d��=�=d�W7��tnL����=�=���\��N%t��o��rM]�7*wq�V��Y�p���#[�uwB�±�rx�{�����
���>��2�6�G=_�4p�l#؜��qQ�JD��N�h�~?�l8�9S�:T��QoB����p�O�Q=�Ow# �D<��$�b|A�֡�&�����*�Ӊ�=]�!P�?k\��ȷ��3��-�Y����o
V��������6%���Pj���V�C&���_��B�� z6����RBO׬��oOO�f���Ro���-�T�X��A����F�E�w#UF h���;��O/ƩǬ�,\�A	y;��UwB:h��<J�+�Sc�~�U��YV�j�݊ڃ(Rs��4ějHqN�Z��B6N�Z�a��2�io.�0h�{�g��K$/���;��sD���;�H�
�l�V���[�����럝6=I�^�d�>Q~�+�����ߗS~�m'GZ�d��(s�M������E�A��Z��{f��BՉ��������Hb��
 ��ZӱA����k�����@��C�{}`5�hb���z�S_�*!
#�A'�d]�8��le�ڶIO�5*ȁK���*.w�wZn� Fw�AK)�F�&a�