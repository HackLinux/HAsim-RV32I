-<Q������[�Y�@���F��eUG*����K�BI�m�Y�i�*[|jr�狫p� ����]�ǁ
�ˎ�$�X>B�)�Yή�*M����7�W��nO��c(���O�g8F��J��*�q$5���`�l*����]a��d� +����L��1��"ҽ����Aif���17��F
h��ߗ�9H���V�]���`/�eQF�z5zv]��ZV~Ӏ�B�\��w��bY���	[�H��Sc��SßsE.���oL�!hbZ+W���v�s��I�*>@�˭��h�(e4῿���z1��C�t�G1�d.o��x�j��H���)�r�� �����5��]ܱ����@�҆���V���v��3����e�|�iu}��x��Ĭ�|\�.β�*��eX�z@�&�����%���MDWz�����{��I�lg�'&5��l�r>�ly�u�KtL@,ր����̓�b�r�%����(�!l!lL:��#$���>�7�V�Q�ߧ �bȳ�=�Py=��ҾaB;����$�2����G��m�v�}�?A&��u?)�ȸl��5 ��I�-�[Ό>S�����P�����?��v|IÈ�&������-���C�L@�C)X�D��;	R��L� �N|�,���o�]��ĞJj�Qᗿx�]��ZaC�-��QeOGtGU_�U�˖�1Ú�y����9�Pei���U_4�JPu�bJ7+7�w:*�����e*{�5��@Dn|��ON5�&���G<�|mߩ�����*c7|�?$�;r�l-�k�����@�z��������>LMe��y]�����s��[����z�t��J�1�1��P��x�eG	%�!�
o�k��xlߔ��z�l�qôeJ�� ���eB����*��A��Jx B��}�&���o6/M�L9�Y)f���sٳm�v�#_7�Ξ�i��J�o@��h2L����v�nlæ����wf&���҃d�@~0�����9�X�ך�.1��|M��0@��E}�9�c%��CaJ���*����n��u�����Z膖o��[{�/�VLF���W0;r�`�r�-Bt�?`�@����Ő�m畕iҭ|"���q��s{����@�r�
o�H|��k�魤&��D�Cf�g��C��<����,(�
�GI��z�>G�De^�ن1�{�n����h%l6�81F�����+���7w�0{�����f@N�L4��N�%�͗����Q(�����1N��(T��+ ������^JmF8���} ��5�M�/>_��OTD�	��bS��ѶF��ϡ�I�R]2�Μg��Rɡ|�A(�&�^	��k5�5eg�����٩yΠJmw�bH�X�R�~/�
��o��	�v�o �)Hݎ�^u&�����-r)�l�ST0%�k/[jɯěcᒸ� ������&�m�ۻ�ř16[AE.⡹���A7���+��^e�x[��eȫ	�j^�*G�n�/j��ʡ�J3d� y������5��%�T
��i�V�F��5ɧ�� ˻EX�/�/����(K��+�A��
������ 4�n��-�t�4%id��˱������ˣ��c�Fy�b ��]���c!�d��v����<Nv��a}ωg���_o�-��2Gj
���������e��(���l�"5�d���l-�	����'>2
�,W�S�����&iSR�ͧ�� ط,��&�x�&`�)vr
w(�K�/������T��B�=Ĕ���-�\{0
���)��xEa�6��}W�/�DG��ϦH��"Ym)W"�����4��t�����,�_��X	h��s�wZ� �d�ɐ0������3�i3�Zln�������-@l�b�J��x���~�o�t@���{v�,���r��h!��zD�z���7��U�=#:��OЭ�7�^�_gf��?�U�!}�?�;��vJ������{׺�9��2��1 17��D�N���l�*�0�I�}φ���g���TÊ��(��p����B;9����D֣��i�W�$�����|�@�]��o�fn�����'U� ����A+���F�����&���3�0�L�7���>�h�HF�s˼�S{�5c$�:eV��U�������~T�K���E���YR����4J��DŜǹ�Y