(()01!70*%7*9.<-=):)3-8-=,=1B*;,)A'2K/;S:Lb:L`)3I%,A4&/HCXm@Rf7I_3CY0?T,:R$/J8(.H (@-0 *>(8L1E[3G[):Q%2M&3L*8P+6M%0C%1E$4P0R$3N$/D"*B*=#0A!+=!*;(5#1$%&(&4".<'7#3&4&
&%7&6�&5(5
�	
'	
HXZIX[J[\N^`RcdUhiWiiXjjYkk[ooZmnYkkZlnZjj\nn]pqass`rr\pp]qq[oq\nn\np]pq`uvbvv� � � � � � �;HU <IV�;HW ;J[�<K\<IZ;J[;K[<JZ:GX7DU5BQ2?L5AO4@N0<H-9E.9D.9B+4?)2=�)1;&.6%/7#-7$,6"*2#,3%.5%/5IIGIJM�LNQ�Q?RS4 <<;777851357!A, 02!$=!(C!'C$D"-R#+K,6R$/N"(H%.M +F%A'G#+K!*G&/N'2S%0M.;X.:X)1Q0'/K$6B%6A"2>!1908#5;$7<!4904)&./$("&!(%-"0<$6B"3:+-,2"1:�"3<"4>"6B%9E#7C'59#*-%*%&#$'1.<0?"3D�/A/>"2> 0: .2&+"(!-/ .6(.*((0!.;$6B#3A .>�!1=&7D*;D)9=&14%01#-3$16+2".4$4815/5 1@&8D%7A';C#7C*6J*7J/?W/@]2B`3@Y/=S0AX6Lb2G^&4J#0A#0=#/=)7G,?V)9S$1B$4B%4?&18-9$6B%8I#9K(;H&7D$5D'8C$6B!1=.4'-%/"0<#4C#5E*;J 1@ -6!+3)7$1B&8H#6G#4E&:D"8>+7 *2(. +:#2A-@M%3C+=O%3E%9E%:E%8E$6B#3;%3;'5=&5B':K(=H&:B+<G,@H+>C'9?#3A#3C(8J)<I*?J%:I(=L'<G!3=(;H%8I&:J$9F#6A!19%;E,?P0@D,6: ','%29/?E,7:&2:#1=0?.<!0;%5E*:@"/4!-1+:%7I+>O,>L+=E+<C-<G/AM):K&:L(;H&7H!'9%0E#+A&>-:U.>X&1Jt��p��p��o��l��m��o��y��w��x���z��v��u��u��v��u��q��s��t��q��p��p��m��k��l��t��x��w��y��z��x��u��v���u��s��r��t��t��p��p��o��l��m��p��d��TnxG`gH`fE^eAZaAY_BX`�A