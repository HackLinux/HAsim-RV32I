300253/(%%"  .DZilml`UI<4%	
  " 	'.9ABA:54372+##!
  ,?R`fhe^RF<3(

"##!	&.:IHD>84234+$" ,;KX`c^XOG=2*$ "#$#
  &.7GEF@;7231+%! !-<HS\\WRJE>5/)$! ###"""'5FGB?=70/.+$ 
 "-:FNUUQKEB=50'"! %,...+& $&&&&%	
")3=C@=;7.,*'#  +6@GKKIFA>=4.$!"%'/8;=>8.(+,..,&! !%'1:<??:3,&$"!   
",4:>>??<84*'#$(09@EIKD935580.( +-.,+27<@=70*"     	"&+/1440)$" !%.8CKNQSMD=?@@<5.'#%'()59:745:?@94-&       	!+'&"  !#*0;GQWYXTNJKKLHA512226;DDDB>@CB?5/)"	           #&+1:DP[a_^XWWXXSMEBD@BDIKKLJIHGB:4.&              	#*.7@MZ`cb^]]^]^ZWVQMNRRNPRRSPF@83+%	                 "&,4>JVadhhddecfea^\\^ZVSSSSSNG?7/+#                   (.8GNYbfhkkkklnkeeed`YSQQNQQKG=6.)                 $.6>JT[aaafehkkmjefc^\UNMJGKKKE>1*"                $+2<IQW\\Y\^abdcdcaZRLIEA@<=BGGA9-"                	 (/29FQWWYVTXVY]]ZYTLD;52.-++2:>@;0$                

		
'05>IPVXRNKNLPRQKH=3,$&.35/#                   '05?GMPMD?@?>B@93)"  !&&                           )29?A?82-.110(#	    
                             
$)041,%"#"
                                        
#$!	                                               
	                                 ����    @   @                                                                                                                                                              	                                                $&&%"        
                                 	 +48>ADFFEA>7/"	                                 	"+4<AELSZ_dedcZRF7$	                            $-.,'/9DGLTUW^ckr|vvrfU@,                         	%/;@FE<3'! !'/<CKNPTVXV\bkty}|vkXE5!                       +8CLOV]ZLD80,-5<?AHKKKJHHMT]fovsoeZH5"	                     '7HPW]ellf\NC9579<<<;><;6679?HVbebe^R?.                      1DT[eiqwzysgZND?;9710.)&$! &-8AJNTUVOE7(                  &8M[doty~���}sg[OH?74,&! &+/9?EJMKC;."                 +?R`mv~�������~qdZMD;3+'!!%&,./,-17AFDC<2&                -EVdtz����������rg]PE;1,),/3555/+)-6>?@<2&              1GXgu{����������|tj\RD93/17;>A?91'$)48980%             3G[ku}�����������|odXM@95357;AED;/'$%,0,(!	              0FZgu}�~|||�������vm_SF>63015<?FE<0& !)$!            0EVenuuqoqsvy{|��|wrcUH?5/++.4;@FC9/$	            0FVbelfb`bfjkoquywusfXL>4+%%&+49>?>7*           "5GW^b_XUPRTW[]`ekqtoeZK</'! ")/7;=7+           	$8GRWUPNHECCEHJNT]diicXK;,!!)/453*

          
$6DMMKE@=851457<DNX]c^VH;+ $)-/* 	
          
%7CGD>81/+&$!"&+4?KT[ZTH<+!$&' 	          ,;CC=4-%" ,8ALPLC8-!!     	
	         '4?A?7)!

'3<EE@6,"     	
        &6?CD=3&    +3971)$            !5AKMG>1$     '-/,'$            ,?LTUM@3$       %((&!	            0ARZ]SA4(	      	 %$%!	               0AS]`UE5+!      
 "$!            

    4DT_bWF8+$      
 %$"            %8GV`bXH;,$      
"% 	           
   +<LZ_bZM>1'                    -@P\bb\N@3(       
             
"  -AS_fe_RA5'	        
	            	
%"  )>O]igbTA4'
         	           
"'$  "7HZde`TD4( 	                        
$(&$  -AS_d^TF7,                            #'(*&"   !5FU^[SF;-!                           $*+)))%   +<JTUND9.!                           &,+)(*+)     .>EHG@8+ 	                          "")//+&%()*"    %3;>><6,                          $"&')*,3.'"!$)'    +14694-                       "',.0/--)" #%    "(.33.)                      	!&1232,)#!	    $).,)$                   $0240.'#    $&&$
  		
	     #130/*#    	 	    !+/-+'!     	   	 (*+)#      
 
 $' "		"" $'&$         			"(),-+&"&),'!')(# $%#	                  '.34530.1465-$ !"!$(01.)#$##	                      $)39===;<=@D@=5440106842,'$$ 
                        $,4=ADDCCDGGMLHG@<<?>8751.)! 
                         %,7?FHKOLNOOUWSONMMHA<8631*$!                         )7@JNNNSSVXZ]\VWWVPH?97430(%"                          '1>KOTOMPPTXZ\ZWWUPLE<84.0-+'$                        	 -;EMRSMKKMOSSUSRKC>;50-'&)*+&#                        
&3@HLPMJHCFJKHHE<5,'""&($                         
!)6>DHEC>=9<?>96-$	 
                            
",39>;3..-,/.'"
                                     %,-,%                                             	!
                                                   
                                                                                                   ����    @   @                                                                                                           	


	
	   	
                  
            !&'*+-./0/.)"	           			
$),.26:=AEGEA<3*						          !#!#),1779>AHOWWXTMB7* 

        %,0330+% #%).279;;@GNW\`b`YPC5$
        
#,28<@DE<5,%!!!").23436<AJSZ`aa\UH7%
        
#,7=CHMPPJ@4+$ #&+++)+-17@KTXZ\XP>- 
	
         $,7@EMRVWWQI>5-&"!#! "'/8@FMPQK>0"		

	        *3=DKRWXYWTPIB:2+(#!#! "%-3:@B@7/$		        -7?FLQVWTTUTSMH@95/-*'#    %)1541)$	     
+8>CJLOQRSUUVTPLD?<83.)%!"!##"! &,,+(       *4:?EGJKOQRUWWUSNKHC?6/)%$%&''%"%&$ 	     	"*08=BDFIIMOSSUVTTRMJE?6-(%$"#&''"
     $).6:@DFFFIKOQRTUUVSQKD:1(# "#'&"
       $(-3:?BA??BEIKMOSWVVVND;1' "%$      $(05<<@<:9;?CEGKOTVWVPF=1'  !			
	      
%,28;=;85246:>@DHMSWTNF<1% 			     
")158:9761.--158<AGMPPKE<0$
     $-48:9841.+'%*,/4:AGIKHD:0$     (19<<841,+&# !&+29@FHFA:2%    !-6=?=83/)'" !)18<AA>81'    &1;@?=7/+'$#)27:<:71)!!""   *8>AC>7/)$"&,03564/)%! "$&)'"
	   /:BEB>6.(# $*.0223/*'#%&(**+%
   #3?FGC=6-'"!%+.1210.,''')**-+&   #2@GIF>7-&!
"%*15510.,))*+,--,%    "0?GJF?4-&
"&,17620/-+,+*+,.)#
    #2?GKG@5,' 
$)/357640-**+*,++&!   	$2?GJH@6-' 	%+2699741+((()))'# 
   $2>EJIB9/)!
%,27::73.*&%%%$%"!	   $2=FKKD<1( 

"*049750,%"! 
  $0;GJKF;2(
!(.2451-&#	  
"-8EKLE;2&&-00/-(#	  )6AHJF;2( %)--+)# 	  $0;EHF=2+ 
#'**)%!   )5AED<3*!
$())&" 	   ".:?@:2+!!&()(&!
    (18861(! "&)*($"!  	    !*021.)  #')*($"

 ! ""    	%*,.+'  $'()&# 
  "#
    	 &()&$ "%%&%! 		
!    "%$" "###!
			
    ! !""		
    !#$#"
    ""&'"    ##%&" "!	  
"%&$%$#! !""!$	   !%&('&%##"$&'%! #"
   	 &''(('&%'()+)&""" #$"    "&()*))('')*),,*(#"#!       &)*+,+*,+,,,-.+&#  !!         
!(-02/--../00/,'%" !!         
$).212.,--/00.("           
$+/021,**+,.,(! 
             
 %+../,*)&(**&!!                %()+(&$" #$#                  #$"	                  
			                    
			

	                       	

                                                           ����    @   @                                                                                                           	



                     	
            !"!$%'&"			            !#%'),059750)#

          
$()+.17>EGIE@83) 
         $')+*'%"(+,.2:@HMRTTQKC7'         %*.258:3.%  %((),38@IOUXZWSI;+        "'.39=BBA;1' !#$#%(-3<EMRVWWRC3&

	         %)05:BGIHF>5*# %+3;AIMOMA3'				        !+058>DHHFB<60*#!(-4;?=7-%       
$.468;?BB<;;862-'$" !!" "*-.+&#     "+12245676799:752-+,,+(%!"$&%!     "&*++---.356:;<:877766/+$ !  	      $&%&'((),-2489;;;<===<80(!     "&%"#$&())+/2778:<>AADB<4*!      	&'$""%'((&(*.2579=BBFHD<4* 
      %%$%%(()&%%(+/249<AEHHE=5+!	      $''(()+)(%#%'+025:?EHGB<5, 
	
	     "(,-,+,,*)&"##(,.38=ADC@<4+ 	
     %,23210.,*'%  %',04;>?@<:2* 		

	     (17:871/.*)#"!%+16;>>;83,"

    	+6:>>:520,*#! &-38:;:62.%	


    	,7>@?<720-(##,2798853.' ""#			   ,8>AB?940+(##+2788642/*%"#&)+.-' 

			   -6>A?=83.+'#%.49:87450+)'*,0124.%
				   .8?@?<82-'$'17<=>:730.++/245881* 		
   *6=@@=80*%*27;AB@:62/./368:<:4*"	    (5=?>=4/(" *28<AEA;75112469;=:2) 
    )5<?@<4,(! ,5<ADEFA<630157:<<72)
		   '3:>@<3.)! ,7?FILJD=71.0379;95/&
	
	   $08=@=7/+#,8AGMNKF>51..134631,#
	

   ".8?B?91(!)3>GLOLF=6.*++-//.,)#	

  *7=B?91($2<EKKKC:0-)&'))*))$ 	
  &3=@=81%#/9CGGF@60+$"##&&&$" 		
  	$09??70(#,7>DDA<4-(#" !"$# 

  *5=>80*!&-4;?>=72,'#!   ! 		
   	%2:=70("!)/6;==930)&# 
	

	    -585.)!$*28<><91-)%"  	    	'/11-'"&039>>;62,'$  ""%%!
	    ")+,*(! (05;=><62,(#!#&&*)&	     %&('%!!(/5:;=95/.)# $%)--)	    !#$""!  '.3778820,'"!#%(//+
    
! !&)/24541.*%"$&*.-(    ##(+/111-+&% !$)/+%
    !!#%)+...,($"#%)+*&	    "!!#$%''+,($" ""&%%)'!	   
!!"$&%&%%%#"! &)))(&%"   $&&$!"   !$+..,)&$"	
   	"&'%$" "%+132/+(#!	    "$&&"  $(/2541,(#

     "$&&$ %)02541-%      	 "&($! $*-122/)#        	 #')(% %(),.-*% 
         #&&%#!"$&''&%""	          	 #%""  "#""##!             !!!""               	
                 	                  		
	
                    			

                            
	                                                      ����    @   @                                                                            		                                 


                       

            


	           
%*((%          
 &,27:63/.(!
        
"$#$
 $,29?DGIHGB8)!        	"$)*,/+&
#+.7?EJOSSQI=."	        	 "%)/3643-#	
#)/8