i!B.]��P�`�Aph
@���q�LD�e��j�݅O�pa�$Ű���s���>`a|%�X� � �$~q�<�����vp*��`\�D �
�<i�tA ��F�>�M�B�&�!��� #�t!�<ǰ�O@E]�`( ��1�Ǝ�J>��CD���P��Z�_$p����Ro�:�H=��2PO��F��R:È��!$ؖV�׉.P�q�����wЙ�*BB��Lge ���(b���=�x�/��ib�"D�n��~Lc/*5�"+�S��,adF�J%�E�aʛ�H�in�=I8�@�(���x/����9�@��r �=8 �3��_^���-Ux2�$?S�~(����R�6��"�w�Q�:�p ����	�����d��/� �"�m���>�9B3�n�bj_�t tCPH�7��� �G���C��,� �o$ؖ��&�`4�  �@]� ��=��|��������VH5�3D�|$�`�H���P;H���emD���:���c(�_Rr�J�8  :��=� ���g�6����P|��D hO
 �&�pR ���Z���>b�E!)(��3���L*�`s|.Ř�C� v f`!�����} >�4�����n��T����B��c��@6������������& h 
`N!" ���@6�L��a��X N`S�����*��A�+� �� a��������A�!r!�` � >��*�Ӧ"$:#*�DD�bX5��#�0��"
6��JdĽ��j25�Z BDZ�F�h�Ʋ6f/�f#�jצT�B�P�Bh�jbԭ�~��E"�a��`� ��H`j��b� a� �at!���yL����m,��v٢�@ �6��"A�Z@ � �Ij��dBp��@.  �>E���t$�F��!�������G:�D50���k&`4��P��@ �^�(
 0�%@@F��\��=#@r����������l!�T�V�X �	`:
`t/�z�&��|��)��]2 f2��(1f�^�G+���JL���%j5hF5� F�/b�v�a����
@@H�*�O�j�OL�K�A�P��%��|!�.���.��
�����X@5��_��Df�Wc�""�A��a|a�Av|��� ~ ���B �@�u'a�!���@`����� ��3A���23&as@a��� �Bl@��!�Y������m ���D$`$>�!���<jn5N^Yc�ec^
BD�Xq'(0O�^rk� �l
0�&�^a
6'��t_�:'�t%���`��+eҾ�Jan�)f�,b&�v4��ة�=�zO�`A$jEfE₥�c ��$�ޤD45��&Bfj��@�.��4�B]h2_��3�D��� ���
�р
� � &� H�1��gbD ��P����  A���!�!��_�n(�J]�&D�/��=I�re�"�����al���Ů@� ����&B&ˁ���aP��A�U� � �
C$a�R�d�E�rF��W1<�����$��A�� @	 �@�
@X�0��{#E�.��!�A��!]�&a�*2V�� ��^eBpA&���@(�aB
j�M^XA+�2i��d��P�,�L� ħHu�  �
A�A�a��D��"n`t`e F  	����v2�E�O��]�H]�T�\m�<im�\`������d�za��D@�` �.��T`J�S ���   @�A����<a�`	 ��
 4A�aX���`�� n� |\��ZB � A�P"�v �  �d�^A�Კ!�"�$� �g��> J�da�a�a��N���a�!�@ V��az��P!�th�O�2��n�Bx&G�D5&�D:FF
]!�us���"zg%F@r"h`b�&�UF��)OTC��]�ϋ�ۂ8abh�E?��Dr�l"a��\`9�� T��� lh�� ��������a�� ���������  H�`S#K�  t�FIb B�$�A��` K%+��B:�y:a� ���a�!�UG0#A�A�a��X`( `R�:@
@> ò  `��3��J*'@HO_#6!�a�A�rx�v��A� 4 ��4	�z�^n+��'�JC��D(YZ*B�����n)cRaFFDdN)Mj_TS
�8���Lg*N a�A�t�`"�.� ���.
*������!x����n���d ( ��� 0 �ybX��r��<CE$���h�V��W�)�	��`�y���� br�(a���a���
@� �
@D�Jtv(r�}bN��6�dkJ3�@7��A���]b @�< B�,�������7��)a�fA�@l�üݓ�i�5CT GDBg��e4D�z^�����)g,��QB �.#1P�BNjҨ_B���e�E�>k/SDJ1y{A� _ƌid/�-�D$C������csV]
�$�pzfW�~��!��DtdC *8� �*\�� ��D� ��@�Kz��-�W�0" ��A������L���,2��# )������(@�t��Q�a���A,�����@ 
 ��t`:� ����`��F������~a�b ��ڛNN�#`5� @��Saۂ��a�P J@�
�T n@�;M+��a�Qm��@:�����a�2��R3�
�I���F���__��%.��$�r�@f�&Yr|A��%{ ����&D��!�aN��!� A˅��@�L �f 2	`��l 4S���H�O�μB\^E�i�$*�ab���a����c�	���-��������2 �` F"����]`~
 O)��xaV��V��`j ����� <a�@�2<k^��| V���Fa�a� j��f�z�υ!���!� �.� B�� ��A�M `�