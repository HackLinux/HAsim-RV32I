�b54�l����4�����<�����V����T�؂%�ivw�'���S���B�v��t���g����HO;�Ot�s�a�XM9�#�i�����istbF���_qfW����o�y��K�?"�C�]8�%��_V��ma�_�A�QǴ�l���n
�(5�6@�����13{�J����aj�jޗ�k/c��b����u�Z�Ϛ�Ū!�#�3�H�-�o���c�4|2���(�n������
�h\r8��ԥXѕ�W�P��>�����P��xI�E|K���T�B��KT�GZ�Kff%g������EJB�U�9��_��qI��V�!B�Y�ma�t♟��f\�0*�O�8ƟZ��Q��q����K�*�QJ����d���2��vB��9��5Yw��:��9L�:3��݋*���z�%N��eR���ʕ��d��l{`~�̩a[�0����K-�IS�����з��{�D!R��iv��^���AZ<@L�>-5�X��F�D-g� ���-���LG!@)*Q:$�е��i~T�9[S��ɏ���F������Q�x*$�Q�� �[�N�>��t���c��2wF:�)��Q!������A�%���$�U��1�턿��Q��d!�Ǻ���6��܏�B�dŦ)�4���(\��mXF�ag|2�<Ѭ���U��&o�po�(T�,�l���hF��HMR75�����4��$4e���������_���'� i�R͈����>�c#f�V߰�$�eKI��tjው*J�������j�nlĆ����fpDn��΀�)�@fS�ݻ�&�L� ���w��}ο
��)'���B��7aj���@���o��҄��5���Q��l�I{�e󤟆�`,�.[��w���ҽ� �p��d�]��u��up�5vl�i���W�t�H�V� ��r�{�RJb.��P|� �ݹÒ��{W �k�?����)6q��ѯ�i�Z���4�M��|o����]�MfR�[���t�xG�m����as& p	�t���lY^���:�iN��&v�%r��&��Z���#a��88��f�#�M�j��6�%z*��pJJ-�:�G-Y��[H���lM)��%�g!A���D1˭�)���<�!�3��.aͬg�f�=��5��3�c��|D��a%Ŵj��bѻ������|��C������|�U�ӳ��K��A�4,��ܩ;�}̤�b`�l��l7&%k���'I���g��Q{5�V]`���$!���!a�E��V`����5��(];��n!�DZ�\�F�s����v�s/ͱ���D(�t6�V��s��k�ҳ-�Md�s ��[k�:�\����.d[����Z\���<ͭ�v�i8�O���n-��y7"�ۨ��[G���PZ����sus��V���pZ�����������[��g�����Z*�f ��� 6�O�&�$����/����!���uˏ�T&���~\
6G��ď-,&��o���V�O��q�{�
���!�4�r����/��eU� ���5���_���R:  #���f��#R���븍֋�oa���h����&���U�d��6yN�g���W�����Z;x�9�q��Ru*������t`��rep�Yek�,�>�M��\��f!#b	�Dd�ձk����zŜ�Q�������U��ڕ��f�N�`ۛ�/2�$�����g�4�գ��5k��At-��G�B�R���@�tr�}����Ř�&T���[{�����9]��d%̘Uۻ�����J���##��)j���b�y#ʏs#ʏ�m��0�b��L�\���A�vD�lqf�Xa����?��������c��J��a����YG1�YnK�͖jo"��٥Բ���uq��l�zd�i�1_V~Ç��^� �NZ���\2C��L�n��¥��|��>+=�3����.���h�J��Z{��j�6h� ���.]jl�~�HV��Kce�@��C��S��Y�`4��C�'7���B�=b��f��d�䆼���Q���P�d�i���{/l��QQE<��:j����������n�&�l���UF��f�^�{��o���-Iv��g�w����t.�+r��M��u�P�5��v�%i�j����kA�jz���R�x*����/���qh�,��vWK��q�������:���*!Dż���&\`)�@�[�r��l(�K����UW�r�D�oc���kp)᥂ص�	���&���r>���
��e��i�[��f'2��a�EY����#ZRs�s��潦���)n;�{���W��g�{����ڀ�:>����nf�yx�7����d�=̠���k����e�:��~oܐ��ӡG�͓���#�"�{3�|ˮ�s!�1�s�E��C%��f~��e���wE����̩�j�g̳�k�f�&��)�X��F@g�+��ySB�+S��!��>�ؐ�3W����Th��1G
�ܔ��X�\���� GH9���!��s�ɂ540{�w�{��Ƹ�1�{{M�u���ǨB���b�d�'��D%h
���%լ����[���Z\��y[��$h2�|������K��a
r��7K��[���n%̘�"��	�O�\Jvg/K+�q�����}��Zt��!]�[����`�r�UQg�#����'�,��Ժ-Qc1X���Lq����$�e<�Y�%Q��
��a����p���#/%��q"#��í��:ǡy6��0В ������>>�d��^�����t$OtԻ�'�W��"7퇣U�ᔨ���8�D��Mr�pב�
Q��2���x�F� ���jBt�[�������l���Z$s�:��*u�ti�',0�g
_���!1�r� �"�Ȃ�s#����
�a����j�qS�7������ ����6r{T�&RDφ�Fb*����R<kQ]�겹�J����X0��
��F\��I��`��/<�� F�Ă�}�<�p�B*���DxJZI�n�,��Ns�G���)��M����h�\����>ұtC	��+&�gA��?d�0UmTY����MUs9�����l�G<�YIwB��6s\��	����z�����������C14����d��C=���}+���Y����iC/ˠ���yx�]�Ԣ�?����s��h�}���H�;�Ĥ�,r�� �+�b�P���`
��D�Ǚj�	���V�0�\��r��1�T��X�%s-��[jb�\�C��3���J�
K�4�ܐ8�
N�P�QW�7*-���r+�k�+���f1d�*��t���׭��t����nX͓s\��{��s�iu�ƭr���v�1�T��~��Q�� ;�Ɲ����%ZF���b������������Q̮���䩾O����oDe�h�"��2�d�?�=��.���]�;Қ�&�a=�f�g��#�xS�eS�ddc�C����_�����r��h|	��T���#����vˮ#K�Cήy�њ�w�/^εD���^1C�fXWvQV瑺,�3��;M�K�*Z����~��'����{g5�HF̬�0엾�����M�ナG�f:��(���JDz���.('�+�<����w�Tjm쿨B��#JV���[�B�������Oj�gʄ���q�1������e��bk�؜σ��+�1���N�V:�nXyH�6��a��$A;�����c��ib��?b���n}���q5�N�ezU#��Yh�W�f^�G�B���4�uA�d@���ob�y�~Nڦ�K����-��g\8�z�[�����CZ�o�>D�����5�y)Wc�|����i�����R��[��Ɔ��)Qus�����]ݛ�"2�l���dǶ�-�K�[wb8��ԉ�q���V�����gc����\c�`���ml����ȗGD�w�����W31㑆����1�
����b��s1�a�pX�B�mu��+Q�%R�*�i!�Z�X��wQ��@t<��C���3�a ���Y`N�f�$f� e�����)����d[rL�4�%����m��`��$���6���Ø�!=�g����k���e�2�`�=��}�'	ˏ�T&�%��2J���%-gS�h��I}Hǋ.*�X�a�ؒ���C�1�n�Kp�7���ܨ��w�{톆+�8�+��
�*��]�|}����wi��3�����]��gE��'�=�!�{}�'MU���,������o�Q��ݯl,�� �m��c�4���G�"q�ᇪ�gUG��^���1�}��-l��e�`/������� ��<p3`R��J���ð���6�Z�P�k�f����������j\#q�Ft�+��`� H�țF]9�q;�v:�w�i����_BIǣg5�K�D�!M�O�!�l�E��:u�&���i{��6�&�u�8��������1l�
u�-�l�g��[��g��x��h�~��%H�関;��R����t��`�0�I���l���r�`����{�y'��}b�.�	a	ƃ�WjüC�p�{�0�ƕ�
U��,�F�c�`Qד�u����_�������}��;��<��W�S�2��/eee�%�b���bX��*�M�J��:@�[�r����Hs��/�_?ƕ�$?$K���d[ �K���ɩ�[�x��#k��C�!�l����`{J���M�ƘkG����ᛤ�����>	'֯�+�a�0o[�whG2�/&uK:�!�2��꧗�s����4m��e��u���L�g
K��<�m3�k�&��W��C�,�`�#���N���`��9GF���<�%�]$�������]���l2��f�~���м�����n�:��%�e���.��d�+�s���LZӥ�r����(���L�c9�t,�rw��"R&����K]��6�c��c1�[b6�8���lp2��R��lBLu�~ƌ䍢�
�!�S�E��g=�����D�RJ�b���;m�S�$�]��}��*%��ʼF�O���H!��R�+�:`�'��C��~!�%0���L��[���`D��BvaX�]��-���i�j@C$�n�f_ ���N�}��}�7�d� [��Y�w��A�Ԅ��7��5p,����s�l����kC��B���>C%\�磧 ��B���r-y����������Z���\m�8��Ue��������x������]Ʊ��rE���Vn5느`']�j#4�Y������R��a���)�Q�RI�L	�Mr�b�y���W�|ò^b� wڜҦ���/�є,�|�P��w��AY�!�E��nSm2���]�Q1l� ���B�b�B)�fb7�[�e6�R\�oG�,����'��g^�-��er�kjtH̭kZ�-��(��-3ab����A��f��u�p�_�_���.�&@�I��F�~�i4$c#�]�����S�y��[�m�ż��LwÀ�"9�)��4&��3���M�f�ꆭ�=��F�R̓2�k�<����E��e��l��!��mT�*Al�����Fu���T�������?�O�x�ϵ�dUi��{����O�Wz�P�_#���점���0e��E�g����o%��4<��4��N���k'>�֧T�����[5�q`���j�iN�%�k�mg�V���d�#h��� O����3���F�L��q����vcYd��v^��$��ŮS� �ϱ� �"�) 7m�`@�k��mٸ$��d3K�Ƿ@H<�ע���Rx���=� ޅ���U��vC�
8�e�٪��v��c�����0�%��{�b��ݫy���|��'��69��G!��A �����Z�8�*����C��W��+Hֆ#|X��]�A���u9ا}��� �����"��hR啹*��cC�0 �ʌ��.�m��j	cJ��5���YQ�ѣ�f�{����x`�%���ba���NL��jL�=�����iD���A��!T�@��D�����j��!���rB�o!8=Sݕ��w#�G�G��p![�~���=8F�J���^m��%h��%�-UЂ�h��R>B�ً���x��r��E[�����8@�R���c�c�{�&ԯ��!���=�Q:�K������T=a�#:�����R�[`C�L��o���ƻ�>FA���L(�~����O�#�N���� ����c���E+�/��uL ֯���]�sFc�lKG���} d�|��c^�;cN�t>�t�=����!C�mө��a��L{�1��,t�iXF_���z(}���QF,gf(xt���?'ÌS�qqr���=��GA�B��q!ΨE8vG"�^��s%����_�p��vv�L؀�ܾ���a��m�Ii f���&S�����b��v����_P<C}��Lbm�<��c�L35�,޸��b�h`�N�7>�FLf\	�얐�a��I�|�M���ίb��g!�XAY%�7�K!���J��(Ҡ�X�!3ܧ�3ܧ�34�4d�4d�4dD˔�1��BL���������y��m��jX�7oc�B~�=�žgP���*z'����Mf�mk�6jns��,]Áe��r�WGS������l��N��n2�����
��D���]�!��$�]��u0�:��6mk�M�I*��u����9�;B�$R�]��M�GU'�-7������8�"%�l��G���h���Y�dn�:������D�cXFP����7E��oy|f��E�C��D��l��2<�h�gQō���u����d�$�a����#�n��D���6�jm��v��-!�mcC����Ack�z�l��
�C�Z�cUV� h�tM�(<��z��l8u1d�����ʣu�n4!{�K2��W��E�E���Ȭ�\H�1���j�\'�^d�if�on�*�rXf���d�Cb�B{.�K�̦�'碄Yܔ�KG P�D�L&V4��	��	Z�h���Ѿac�ۗ��e���ӱ~�i�� ���5�'ٿ'�!t�����_���)��'"�!�ʢ�9��	:�G[��M�eX��ݜ��u��%@��do�R�f۔��*W%�7j�W^Gl?₏Da�&��W5��f��c���6?sp�G����m��FB�����on]���s˭Rۖ��e���ڑm�<F+�oe���W���,��5gT��r�r������Y$�ӯqE��_Ǫ_f�:��HF��;���5U���^G�!�b��ra󤓖�� /�
�����Tt��<���Y������=a\S���m��0#d��2��rny���6��&C����Z�������c|�Q1��t�撞��
��o��twA;m ���t�Sf����Kn�
�2pg-�k�@g6�Z���ғ�]�)������:��eS��'�U�U$k8����2�>�ՊO�`۫��r�3�]�i�?#�S��lc�N�7�����b�#I��޻��R�P����khc=Z����*s��c�vN�ez`r�oMr��Ϲ�&��aQ��`rJ�H��O�i6j� �ܦ�fm�E*l$�!��tx�ނ�Be�U�����r�$���Ax�a�f�ic�B)C��Q��`�0���x,G�����:�=X#���G��3 �_��v"^Dԏz���ز�Zs��'��'�3���$^���J&��W��zf���@��9%p`�)+e����q�<��_�09�RU�=����{��eC��d�M��b����ν������b��N��几��b�`��d�3�xj0ou���(��m*�}@Mc#C(^v��.Ą�X�D�xrhY�������fS��F��+[p��[Eԩv�|��^�o�leĶ^ru;A�N��B�p���-�[�e���gF:����c��糮��e<���:�
����n���"���0KEA{��Nm�W6j�{.F��&G���Ě8H�5�<���e�G���W�{��$"&L���ٮ�M�KϏ�WҥQD� ;��@Xa����%ME���v�G������y��X�*�����&�af�m�ԏ���̤���k�y?T4���A:�Js}�$��P�d�L��m��x3�2�E��z5Sng����tZ�ҋ����m�_���2�u�����8�]��;����bt�g��(c��_�G������u�b�C>�f��+	����t�hmk��o%�_�W�3������l���lo�I�yʱ�9tK�[���4l�n�	��������p�k~��g��k�
���kD;˶7�6O�n��s�@�l?s�X�"9��^C��L ��(�c�
��ҟȸ��~
痩մ[����^���sA�Uȅ�����b�#���ʖk�F4��3k����u`�m�PD�gୡYЪ��b���(:s�X��8*���nWU�i�A<ܣ��`��YuF�T�	%����������T'��%�+w`��y����tCt� ��P�(B8�K^��9ń/��QȣL��Ǝƶ��?��}��7���Adf�F�����R�a��v�֦�&Gz��$�Q��oC���X�-n*��Uj���~�<Ӊ^���u~@�[���a�� �*��+[Ck��hʲ�_�X��f��Q��G>����!e46ݭ��a���M0��B7�]��`k6�,����C<�3F���t2�m�;_��M�/�¢lz�j0y���i#'H�lo��T�{�9$�C��X� 2�jJ��I*�I%��6"�X
�x�x���H7~���=��-z��n��g`R���d#�_���elL���w�@�FT�����[����rG�_��=A�^�Es=��O�]3�k�5E��L�G���Qe�R�x�yk9�S�?ߐ ��S
{�6�7z�s�˒��[+g�y+%5�r��8%�R���'vJ���] 	c3��M��3��QqX�P���wq��ݿ�1%(�惡G�����p�`� j��B��Z���������G�����������7˦�B��I�\��J�2(�2%��z�Y�#9G�h��c��c��QmSP�������7L#�N,�G�ۃp	c$�9���ߞq^�`�N�av�V1%Zs��H��H2	��M�E6˦�q���a�A�%8r�+��0��%�qI�+;�zt<��X��e��E��s![�[�K�!1t^�Z�G�_�@�7U|k6@LY%]2�N�E�~=���OE�4�Bu4-SL�����k�l~�8�̸h����e�/0lF
u��_�<���$q��������=�RF�'�j��kz��t�a�~�F�sjU�bj��]�<'�`Id���q���%�(��ը���곾'$��fR�����v����^��k�`̵�m��I��� �d�|��5��?�u���*�(��=��-Π&P��ٗ��`K�)u��L�	�@$k����s���yvb����݌�����d�B<'��|�~��eC���î�λX��kB��� H���* ���	��,gj��a�gZ�9$s �x���D�J��+���s^�B������?f�zk��Bq� ����2��e��1kgt4��I^g�U����s �����|f��5}0��״:GF��\����5l��*ݍ=��:��L9:�F�᱃�D�Q����Z�[b��8�"������G��Ǿ��O�=�Y�b��S��:��\�^�b���C��e����5Q�h �uwE�F������,��ԫ�9~&F�1��⳶pF�	����w/����l�O消�g���K���)��F:��t��l�?�4aȥ��-�������XT�ac9�wP����*�Ʒ�Őh��'���7�l��!&���Ӵ��Q��X�NÓ���L�T���8�~w X�]�<�м�$���!�*�f�B�`Ǐ9�#����ww*��o��X�w޾a�@�;�&=R����$�\��67��
X��|I�O���<�hR
��e�5�w�2�]�2��a���A-����ܗ���_�R�!�v��b���̨h�� �`hD�t�,��r��WR]���	��NJ�P��n-�l�}�`�s���a��g�̿�����9m��efˢ��3�<u C6���V�`4��*d�o2����#_�2����b1y%�.l���u�[ǃ��Z��|����	���>�%�C�3�Ca��+av4fD�������Y�t���q��d�خ���_"U�l�����m`�X|�9)v��q���aI���!x���o�E���95�gs��`��������_`�$��8[�,8ch�y���A�|���%�	�������}C ke����|���,��jV�/ƍG��f���j�K����(b����"1t�.�^��ħf��I�S]��z�����U]�ʬh�������9l��VL��5�h!uf�%�j��[�$h:ʜ�;�%i˻�a�e�2�`�=����jG��n	̴Zn��6���N����t��ta'=�䣸�B�[a�e3�h�#�7s;�X����ￒ^��M������5d��I^��`�e�s�������e[��D�1��<���F�N��r,&�`s�I����x�ɚ��h���ϖB�o��pm�������Z��-BR����͡���i ��˘���cDsQƹ�����������������l#Cn!���G�#��sc��B��h�)`V��#���:���,��H�9C_�������H���\�f�~���7j�O��B\��21�2�1l�L��8��P�|�-j��z`%��jf��Z�C{.��I�C���kCݖ����z�&�kq�a�Lj��(�Z~ED'���$2(^�2������5�gl�&_&�j��[�0�pK��=ƥ'�@k�㶧	�k�g#k�$���d��s�����-�0%d��t��g�y�	��Fk5���6�z��c<uB���Zy�2r%X#�5�K�ee�eeY��lhG���t��G�\$�'9�l�y��j��\�!��!�����M��$�����ƅ��q�6ӹ^�'Wa3�䴖�~�s�J-�߬��H��T�\��#Ӫ�'�U�N�J��5�Mu�ͧ�B��sa��ަ��xC
�C��6���{@��;��$be�m��!��ߚ���͕r��`��ia�,YA�,��եs?%Y���x��i�����75��G?tЫ���V�]�����J�5ݿH� X�{��w
��+�jXË��"=�1�S���)��j����"�]�g[,��)����782��+��!F��!�t�nd��� 3�hfLP"�l��ƐlŎ��-@v ��h���amk�!��������&��'���Y�Gxd���������bK 
D��t�f�{�䣂e��;^GC_d��c,����!5������4���{�0�{h���.2B������؄.��a��xF����`͋�i����IY�Dr�	z@�Y_�`3(I"N�����<��f���,����w����li���d���BE�vF��	o��{f�D�Ƨ���v�����u�����.a�s�o��Yi�쉪x�[���{H�k�%�H���s��8C
�udI��`B ��s��{;�� Ef�T�F��Pf��w�����A�:�#��2U��������ܞ 4�����.��ՃS)��P2���/��(畚���|�����*����Z����@r��3#Ցm$r}��:l���+�QŲ�d���� 
^����`%���0�����]^@��$~f����a��'��$[��@�e�c3�X�"�샎����S��Ӿ�c�<��j����X�]�b<�v�B��X*3������cW��W�|�촙�EKg?z���'M�]��r����[j�葦ŴA���%�G,]��������B��� ��_����!�11�	�C�\b���$�C��������9d��o"�zT�����`����ճ�������fֳ��;	�Ƃ]�ƂMִ�����l�r�f�g��D�?��i�e2 r`o�d��e7��~�!������7��gO���R0�#"3��
�&Ʌ���c:u|�c=�������.�u�f�퀀����&z�!��"b������Ws�#8�X��ʯF�m
�@��$j���&�����%�e�%����$����#}%��O�-f�DE�d�檷���
n!��ф�ǖ��ǖ������I�ZCF]���р���C�1����E�1�/����+dH�� �f˝�C�zY �z��J�y�/'��{ؤ*�J��-��$�Z�'�J�:�
4�l^�4�sdM��44��"����&�"��aq��s�L�1�~�bM��eM�j�R�d��ͩ���i��#��)&<˦�"����ᤴ����鵣�������fٮ�lu0��G�<��]������C7������{�㲶ePR1�;4�z�ۯ`!j3���t�c�t��L��懡ES�P�Q�W�k$4��`B����3��ޢ1Ց<F��o��c
����8��6�$�f����w�œ�e!J2���Ftφ22��D�`��@�r��2ɭh��'Xl�䚉��,��l�Ԕ�іf���mI
���	�i�~���M�T?̆���G��@��Aw`Nw�}�iI��`�������.�F.�C�֏��x�䧔����S���VgS5���>S�$U=���l�C�o�c���c4��Cy�[�����2�+�33��^��d7�d�c�d�cL��������"cZʳ<c�	��4�fEN�aK��^s�� �m�9u�z�����Q�#@�~`�~��L��.�'a[����1l�̋��赑��w���;�EZ��M��c�}��p���)�'{(�Oo��O� �"	�W��Oޡi���Y�p�d���a�p�`[��`[�k
�_oJj��5m�Y��e��\��Ŕ>�:�xǌ�TC��k�k59��]LD�#���bFВô7�c[����h��!��H�<F��ha��+Ŧo�M�:���x��,�������,���\��r׸���\� �i�r�]f�ߪ���I��^��-�lTu�(��,q���sc��^���	�� �"���!�m�!s���^��X�l�:(�O�>�R�ƛk'�/ސ2k�����0��Y�s	�qK�	*���Z�A��aƠ��O��1��e��͠��n��D�>dgSB�cd�3Xc�C��m?daŉ���k�hD�x��f8�� ߥ��ʥJ4�l^�2��V{����:H��3T3qb]�P_�I�kǗ��Ϙ��x�K.T�)Tj�&7�(�J�N-�܈8�q�B�R�l�u�����#�"Z�d����e����~�⎉'��W�6ܸ�Ecg�-�� X���hG�e�l�&d�ک�9��2�XE����d���h��)e�o:m��x�RrQ1s}����ڹg#C�H��b@�$º�'������G���k��;�'������i�o�� �	���-��m�k�ȿ���2���H������稍�����9Q����-�O����e��u�"���ɜT������jgߋ�,���RH����d.U�pd��e���E2o�G�s��)P�<~��U��S��-D�'ke#�W�E��^�گ���G�a��X%�����h�nj��&��(%��n�_���T�a�k�U�Ag�B�6"��t=@�NL9b�eX���]��#�����uv���筏�rd�Ԝ<䳈���xMl�i��d���%�1��Mփ�I�#]�����J�s�ڨV�J�h�[D�#1S�Ό�avᨴ
�`���I^�Pb`�|c����3@��qp�k$�#G��T�Ԭ����X!;���t�,D?a�@u�h�A��G���'�֭ک,vON���v;����2B'�7��>�aƍS��2����4T���YF���*�zD�����v���1L��MpFH*Y�F���!�ԛGa�q�\��=׆iw>`������t�ĂI�(gf#��#9
�ſ��'8���NC$��N͓�'N���U���s�rnA�?�B�{� ��9+E�Tɾ��� '�C%�A93�k3c'��:���ʶz�ޗ1@kƒ��V���Tl��l�˗j����W�eK�yC�.]���г.8`	l�Y�g���q�R/�ࠦ\c��t~m��"�<�kׅ0�E�~tbѳ!�lЉ��D�Dko���߫�ʺ��8�nb>��g� �7ʾ�٢���Tf}g{sTc���� ���nR��6k@��m��g�t�� <��5��_a�k���!��L�5�%Ka	�k���tg��٢�3�a@�E@���ۄ|,�2�_������}�Fv�6�Ze����-7m����������R
���%��!�z�\4�V��ѢO+d���y;�3J��S{���T��1�L[ ��&��ӂ9�N$^rR%�q@g�t�d�s�c���ׄLZ�vM�~��Vn��w.�΅1̢6�T8`Na݃n��tE.�Ҟ({��)/|��.����7�-�y��w�'��o`�-N����v�"�-y�+r0(��^��ZKY�d�[�w��SZ�4��}�;�t�?h��FI�����k%m�nj��.��u�+��N{�T�M���*�+��]i;P�������s��pk\T���A'�վ�,S�Ӹ��W�k���`d��^��0� ��vf��fp�m��y��+��5�����j�x�`�$�낖\���&�Ft��;��)���E&��tα�ˌ��� 8�t��+V��I��49.�#�iXH-7�!��4,bWf`D8�D����Fx������n�����f��Ed>�T�g�[��#������2*��֌t�y�f'.��֕����-ʹɓ��j��r����*�������&����^昪�ک8�'d�fǧPb&p�;4��[�ߒ���[}��rv�DrC�xrm@����<uě���5�<h]b4�_趴|m�����ɯY!�T �6יfToCѶ-�L9o'T����F��(=<U#�#��e>BKE��r������L lb�Z�[Z����`@�ϒ�O�@��ź��B�t�h\��,/ጨ����Eo��H
��i�����V�.çU�VB7�!{P}ߓ>e򃪔�T�rz	���<ܽ�[�XP~�*�+��~�pl��b�&&�z��H��*�۹tC���m���L;�ě�7�Y�>#�!<��}Y���m9~N�'zg�& ������n�+�-2�����n���c�y֔ͭ�85�+���+��,�����s���Z�[�C��%lR�p�<p��>.�H{��x��t�z���(>��0Rx1�
bJ�4�Ь�2��*]��ZK�_!������ߕa��翌�3�u}�My�Y(�r{uw��[k9���`;<��c,��ZI��K\�;�B<6]5��Л�u�^�6���7�A��?%�@!r�d:�������|�y������V&��(�$�i~�$��}�
���o�f-Lb�X��}�cy�s'T�������4�4�9���a��F��*�w�]�fd_�nR����#[��Pf�bp�1I�\�
s�'��.t�|g����eUT]��)�˸���M��'(��5�]��Ÿ���:o�o̸�%�S!r榳Q�'�v��c &T���]�W�)�*���U.���eDA_Hm~������b��Ps��-.r�� ��3fK���ʪRЪ|�[C�5�Kp)�	˖O/�aDW'�5׃�������"$������2�ص��!I� GLܷ�����B=����|G�e�M����i���4�-���'������{<_p���9^�ƥ��YS)����``��>�YϨ�#X��^-�'Ec��Zt��%�����i��O�pN5 ?t�b�$��E���#��?�U�Q8��.*e�N3�EN��kW�g_�}nx������.�㹀�xn�G����i�A��A�TG��Xե��7=k��g-bl��Ņ�l�Ԍ�Z����y��C��zy��L�����M�m���������ja���c��(%Y��A�-A#Lϯ����[���a]w�E��
Q����1�����#Ԯz��3������Y��!U�g���C�N7JO��3%��Zs!a�T�j�g&�!F�o�3#v5	KN��;Z*�����a��A�-S���ȁ=7|�V��*�Ǔd}q�yk������'�k�����>�<;��.+bYw`��!��X�|��`��n�s��/��v�wd�Ǡ����g���Y�����Kf�[��pL��.��n�!'�{-�����Σ(�k�#�s5X�bZX���f��g���u|U�م[*ˊ�m� ��{cB_3��R�jJ���y4��ޝ�M],i�;'�Fu�(�����RJ�\#�n0����@2���y�B�i�3��	L��jg�V ��%�>���g𧭴����h�yڂ�{ϼ�}E ��zF߿�����Y!`#;�\3��;�G5&Eo��4B%Ga��Ĕ���哖`�nCW�T���m�'�[�5��|K/���;�w��%�'K����AC%2���e��p^N�������+��j��P�c-2n�6����h������o�_�@�%����8��u�Y���e�di?��� �?삥ѿ}=�p�6�%��m�$�(��o�݈�+i��k������`��D��o��ܰhb߃��c�`����u�jdj�������q`�b��A���a�W��Gg�s�`�n~�4U��+ݥ��ُ_16i�����諌�cy�}1#<̄�RR�{1���(V�s�&R��������2�&x��� �����Ӎ����ng�v����0D8���11�����G&*����X	��8�$!L��{��WG�²H�@�ml���DoF]��垈%����#���+�u�"1������A���]����8.P�P>7!�l,��@
�he���V~e��Q�����M�}m0R�����x;����	E����s񯊣o(���t�/�'J��B:��uN�jcX�2���٣]��A;�L��v|G�ίp���iTb4�>i4�>�x���ɟ��KtT��ȕ�PQ�?�sv�w#���(�K�����:�xJ�R��wɯ��5kk��{1��ׄ�Y�$;�*�T�?"L\��o�Zr�
��nS�e����:V1-���Tx2A�y�	Ļ�pAx�ᙡ�&|.y�\;̚���r$�*D���	~���yQ��P��'خ艭��Y��.����!0��e=���{WPᗼ�	P�0KI/���jk{7A�����p�7���h� ����zN��h�ze�#��
����<�[��]"YZGZN�AaD�˕`�X����zq�7�$��J�H˔�{/7���'jJ5��-�s+�k��鋟� ���u젵5f�~da�	��6��5ȗ�g�8�m{�?����>�`?؋�d��#4�nsE�\�xc��{����`�։$#�b�~���j� �~ɕ�8���x�0����t�	����Q�j����EJ7ݣ��z�ͫ�:��p�l������V���JeC}�����}n��<F`���t�
�r� ��q�`S�)�쯨K�\��#5��^���@�i5Y�~���W@:�P���ŕ4 ǝ_�q�?/Q�E*;}���d���h}F�y���z�=�a#A��B\�d����L�_�wI���!��M<Ӫ��c��yz���B�-�˖��f{��� �M�ӿ�7�F��F6��:��Hb��I�`��l�|�B��(�DrDs�� �Zi�2Y�ِ6D��5lY��/����uj
i��,�j��)�@�9�ZB�>���ϤJ�3d�f�.�@LP�{fa�:�T�����o��"�����d����xI���4���~��.����W't��D����e�e�'�'���pe�ZWc�s�-g�/u�����\6��duC�w����H��j�>���V�����R�	Ĳ�~J3�l/���6[�J�Y&P1��U�3�����0�a9�j
cŻ���Z��Mά����X�H𞧔�ʭ�f?2纈h&�t�*�ku�^깋&��x��S��S��9@q��������?#R��kM�;�G�H�iX��=�����C�o�{�t ��=�޷��K�y�@R�.�խ��\�s�v��"�qƏ&��C�"ƞ�{ԩF��-�
��M�h�~Z��P2�*3?�#8f�˵�ʭd��oc���h�Gf#�qH�1�������nAk�Q2l��e�b�O������_44n8��l8���Wce'�(�a0ٮ���HE���}��3�Q���LQ�d4"oq��H��]����'eO�a[�F���q�����@��u77���A��'A_e�b���)e�L����`h��i�.A��ۢh�"�|臊ٹ�1���j�����b�d������e����l�����Ϥ�F���ŷ�$4#��W�+����� ��j,����Vn���s1m��ǰ��4'C�{�=����R� �m����O��9@Q� X���\�J��0�7�����~���~����fةC�k�v��'$#l����ʑ�漦�1��)���K2`�c��=�{�U7��f�`����j����+�nZ#��\����c� �ل#�wg�5͇0d�e�D ��y��	�w4�/�#�ƊG�ױB�����J�ni�<4�m�y:g{0���'_���.�����X�ﻬ�Y�V��t���w��%�5@������~;k�2����[�`f�t�J��i2��%���xY�l&G;(
���L�aC�Δ�-�Ufdq6��x��[)��lm�c�@ؐι�U��LE�\�؋���4�j6
'��	-�e�i�?��M��X�z���|�{,+ơݥ\�����?e5���K�=rY����T�X"�F$��Fi�h�f1<HS_s�o��Vlt�F��$�ABB;���RV�����j 0$i`<L�"#m�yC?��O�P-�o�R�R4�8������P���ؖ\�H��e#���D �R�EȪ�a���B�u᳊� &o��v-3���@<F���_ ��|d*j��dsGv��L#+��9�t#�Ow��X-�����]���]�"�����P��j��k�->ؿ���o�h�gb�'��[�}��l/�(N�~��L#G�-�Ck5��fU
�D&��XiZP#h� �`Y&9'����8�m�ƦG�t����\�ն�T�&&
����%.��F^��@BEtW�+l��r��d���G�|@�n�!6n�E�+�x]M����PԒ%sa1�B���\�~�ij�|*;�9���@̧
��3usu�n�����B*����N�m��_���*Ct�ʣ��扊l~\�/���Һfg]v<�r��T��������F��!��PS��F� �?cR�i �M��C��v�Ye��^ K���#*`Ĝ��0��S��xӭ�I;�'��i���!r~�����c��,b%�h &���_��A�Z�Z�Y�
k���k]��1��ū�&����C#�7y'�����&�ws*�"G��H%�^,͘��]'<���y����?�u�����OE���a�����3��s�����i��&����VJ�⿢4͟	$��I�Y���Y�%�l`�B���Y��FsB\��T��hj�B��H�$�|�oL�B��St�@�A����)�
�I��ǻ2�͎������� ��6`�%�+�$�/S�D�
�/�&ej= )�s��T���6����Os��2x`9�v���������X�jr.-���Lףj�Y�/3��y�� 3-&w��|q�����kM�3�cg� �*��GZ:	��R�/�bǐ� <f�"�^Q�w �m���p8>�z��à�㗩JE�ei�ʩ���@D?Յd/y�,��4�L`,��u�g�g���T�5�fo����ɌL`�����]� ,;�(<���l<����2���:�ea/����_�jcI�'[d%�Mq��*K%]��;��r����2���֐�e�N�ƘkG�6eB�����"�;�.hhD�+�LJ�r�g�/�N�B����o;GݦO�qY��m����2�ZPǕ�'�Ǣh%b<�r�5Ed+G1�Dbo�h��nsGE׌���ks�!�P�ri�р�Xmj�	.��Ƃ��@amU2�d~���gv�"��:�e�%e�DI������DªiYVox��
�q �g�fey̦��Y[�U���P6{����v���a�ڧ�o���m������w����Tx�8HzZPw�co���,n>mC�"-�3��S�%�qe��N��a��^J���M��	�T�&>�/J#�i(������H�-�q`I;��A���؍��3��'g���VB���c����\���C���;̘�ȸ�����DĜ�qp��Ԁ��3`Y�I3�e3���r���_��_����4�W3�G%���7���_���L�J�$f��ɢ4��BM���B��;G��[�\5�m9��"�+��e�@�0�I�Q9��l�2l����0�2�:�G��X�c�P]$Pu���p�'%��~��a�����'��n�0��m��a�l�ץ	���>�`3��g�!:��;�� >�PJ�	ǰ�,�a�,	��:���qZ��j��	���J��O��
�C�Q9���]�Kr�K!猹<F����7jR�H�.-��Ф��d��jp	�D��N�m=�t�o�_�����XíE9˝�+�l���r&�Ɛn#��J��Y���X��Lr��b}��J��Ra�b�T��@��#�$Z�#��쪕�C ��d���]�dA���~)�0MS
ҕ?#�J,e�<:+?�ZiU��9���S��rc� ���t��~C���=�ƶ�9tK�ƕk	�����7��?A�l������aZ�a�Ɗ��t��������5�A췟C�|!k:��&ʢ� ���'��a�i��������\�.�������;� ��#rL�]�%��������jU��棵#��gj�#V�G�o����$��|�Z���0�L�'�Jb1���P��@t��d����d��Xmí� :>��f��]�����W�e�E�:�����F�#�͞�.ܥ=�ó��m���	��L�u�b��ـB2�5��/�	���%�v�T|� {m%$�l.���4d\��T� I����>��^*�o��-���B�_�Gus%���ר,.G��3u����}9k�ܩ�������f��Q��Ϛ��'��GzY���u�n�2߂���~ct�-�d�&���z�����إ� %��bjo����%l�3Kb��s`�d��)�z� ��.B_���)l�0n�jFx\���A��S����v���R�QY`�Ӽ���(̥c��Ɠ���g2#����*w�x�	�$t%c����Y�����:��:ӄkE�P�L~�qM+Y�s�qJ�]3)3���8�����U�R��{�)�s�k��Uy6�þ?1G�
S����=e!|�T����O�U��� <�oi��d��gz���c����Uʠ�U����zMr�ؖhӜ�'��_���=�z�J��Rx�x������ɤ'���?!)uqqq8 ���4��K}7z��;����D��x�D�sC~���-��z�uݽA%J�g%�D&\T]n� �+�2��r��k�d�Ҁc�����@.������}��Z��o'���%Ċ���(u	�|�R�m. �=�2�9s�rl;�!fZ�e�!qf�zC�W=gR��l��j��DfR@���)%���?z���4�п5�
jT��sb��W��'��}
�]���D2�6���k�c����Ř�Iy�F��òZa��j��M���`W�U�����7��0�p���ussòL���j�o�r����B�u��FJkd��ud���瘿�D�b�\E�&Ӧ�%}�˻���!�
�2��x����[��i8�O���n-��!�Co�?[�������Z��皝P�zl������pZ���o���Z�S�`D*�6�i���������C���ݦ��k����3�� ���,�p�j�tg8���l$�[��|ڸ�Y�\�����������`��WX'���n�e#������� F��d�;��]e�u�T��S[�Ϛ�����\
�g3K;�/[�G,E�58�]��3	飓�c��ͧnw�@�K),�vD����e��p�D�OΖx����j�o=��T	�+�,-I�F�NѦC���	65D'����5z��$��� ���:�p��b8ʾ\����v9��T%�Ֆ[a�n�&����j�Qg�3�� �8ͧ[����\B!�G���\pZ<�o
M!��]��7�2�-m�m��Q��hd��7�wp�F�4���g�xe���R�9<�W���q�r2�|#��|J�~3�����#HZd���������{�@$�bh��wS��JR�^v瀍�S�����H�2���,qf�U�����Ț�>��	����r�����M���i���(6�O3�ћԺ2ȤI�%����� ��k����=5̲M�rt����c��b��V�4�c�!�[��L���W���eb#�	�>�&���$����a���4��%��x�y͢�@`y��z��@L�!�taOlh�%j՚)揊�����bQ��2��5�0�o���#��J��� ����׿$!�} ^�b��c��a>�s������6����m�`'�B���@>Č�����
�d5o�����B��Yc��C�f�2��������wd�t�aj���e����U�Ʌ��a��3��KꞳ�D����q��G=���eޣ����L�"��3�U�B���ck�)f����,� ���˃DK[#eM�����2w����Ξ���A�S/EhB���[����@��º`�h���=�"��m��Hx�Go�i�2�ɣ!0��c��Q�V��.�:,�Q���_����:�!� j��у�a��ZnD����lz��¸`L+��輪��/ׂ�Pbc�eQ��)�ρ�̃Ɔ�+�i���$'5FM�ny����x�f���O1�Mϳ�uq�tF���.�3�G����a���=�`�)H�)0�N�P��ecfOhGЎ/��������=d֧�A�J�vHϼ��Q���ὶ;x�����P��J)P�8O��@@��(���A��C�k�v'c���IVMB��N�sn�F�h�� �������NQ����̇
��ǣ%92�f�h�K���N`�\�J�/�ro8 �D�D�NĤ��qU^7����+�QlN������DF��C�MVΠ�mIVwh�o=[-SD����ED���+삈.8vq�g3��;¡�^�̹b�͹b��v�ėE� ����pX`����l-͍7�2I[�S�t�_�m�i��B�6S�hQ3�����q0��RD,��d�`����g�i.+#DZd�@:f��ǲ�fYs�F��I�-�0�"���"����K���b���y�GC��%K�i?���d�J�j?���x|R��!���mب篋&����y�U�g��Y�>����_u�HD��r�m�(�.��S���#�͢oEci��������f�c����x�ͧlc]�0L�ݕn罡"������"��k�����t�%j���
�m�dy]V�|���c
P��5�4��\%����<��D�TƖԒ�X�-��h��Wd1��WcFRW��ʊ���c�d�e�MS���)�|+����Tc�Ԩ�Q�6��/�ZإG��Ǜ�g3q���������c�o[�]6�4.*��R�-B�*Oa}��L"��8�-����aI��by��s�����U��e`C"#3����
ŵ
���1�0�FD#����R��"��z�FN�ub����A�ܶK������E��>?�&�Dzc��bǼk�٪��ǁ$��,������%����^�"��#h��#��c�Լ���%��Z�]�B�BPb�[*�ȫc"�#n����}o����wᾥ��9�B���B����¢�ē[��#㫤Rć<j�����3ʊ$x������>��N�\���k�{�����Zb�|��p���C}��.�c
�gJ�--ȱsB����}��Pſ��v?�Dέ��.�u�na��4w��h�������re�D����*a��$��-��������cM"#�%̕C��8<�Ҕԣ�e�e���>Խf^�O��Ė��[�'����wSm��t��?��Q����6�$��x�'�h�wB��f�f��ϥ�b=Q�%P�ʾ���fS��Z����]��T��C+��h�;���P��L��ͭD������('��"c��B���i&�))��ƌ�d;W�;Vb����ٸ��`#���g�b��>Q�8W�:��s�����e�������b)b��d��t��j'�k�jb_Hm�/@�����dp����s�+��eְ���t��x�h��G��ݫ�&��8�̀���G+w�n��H[!�U�FE�����i�'��j��+5��3%o!���ʀ�o��l���,idt��x���&Y�\�)۲�8�Q�j�`��,ݦE���;	�U�bDu����aq�6�!�6�d�&�gـ�,����,䮡������BZ�B<F�	���m�;���Z�;kC�#Ŭ�����ỵu�����d�ͅ5�"�����<�f 6ED� �@��c!���fbI���ëݦ����㵚&P-�PmlG����Sآg��\X�o��m_ĥ&�J����ݣ��M�