�����'���������<��#�a�����geο����y��G�B����l����l����z��3�����şR�{�K�ӝ}����ˡ~��0�����U���O��w�������iEi�yU;tj%v%�����'��2�|֡(������L�w�q9�bBi�@p�H5��$l���/��w��b�v)���_J�Ǉ �M>�}�����O����o/���������N�-�NG3�qv��B+A�ƥղw��"���������y�3����������κO_�W��v�C�L�����*�9�%H(.�8`&(�GHN�U�9���PDN�0ɟ5��a�=V��X�"\O�Y��ؔz�pLPK�Ny5pmY���#�����|�y��0�;�9|눟�~��IJ53�5k#�2늎{��s�y��!?h�N�T��Z6����0��L	M��
|�S�Y�I����<���$�����a�)�h�d3|`����tK\�nSaj ��Ji��I}�P��	8KK� �	rTb �t����MVYT6�T��lp&���9�jhC@�Mw����9EM*W����7�-O�R{��YÌ�m�>��f�+b8*O�o�x�V%�O��8y��o,�|V�\���]H���Z;�z[i��NJ,Nl�S�ҥ������~bEv��|�c �	�r��6�׸�X(D=�O�t����>φ:ۓ�+�+fOҶMǽ��?tq�)�)@��#�\M>�Q*~�Zq������#{��SpO

��'�rx�����'73]�����3)��L��i/-v���n�o����c��� -�5���^�'�A��6��`�_���z	��(a��=��9�$ЎPM8��D������r�e�L�T"�2K&�b�bx
q��ei�"_wO:>޿=��x�4�~���-���^>��Mx��,���ߟ�����zS���(*eו/�v���V��ZX���<�7�j�����栗�� 0���Ʋ+8���|�ui�c����r�Bs/��V���{���L��Z�\6�[jO�@�����M]7[���
�~�Wl
��
�9��x��<���?�������ĪW�������4�ސMH7�����$�^k�v>��S^�i��%he=椪Vͻ?Ui�.)�vx��xO�|GFY6����|�,.���/K��%��-5��N|)Efo���u]9G����E��
�o�0�ݑ�_���5�Dd��
���������Z�5slgl/��yڝ���e=����)�z3���mh�����}c���]'��W����JI�I���j��f��nܘ�(���{�)�*��~u;?�.ث����s}y�6�1ā�t����S��"�E�h5��U����zz<�:�ν���=_��+V�V{$&ԁkLyr�xus�mt�3vY�kG�E�m�-Y㏙��"�(��R^�-�~��C�O����!����Jf�DZw/z�`cI{��H��������*"$������~)ԧ�Vʜ���]����E�������X2�@l̊�>�������qg���R�NL���s��=��{S�Ks�R�ڽ��ڕ����m�B����?]��d�=]�]u�4��n�p��u}�<I�hY>B�<�kW��㝢�*^����ΎvsJh0)���r�|��{�9U=inlNm�J�z���fx{�i]-\+�GZ�ri�֊��⋝��u���(N��PI�h��)=�{���5N�2G�*�ݘA|�)i�^A<�E���rSӌ���z�3m�⤧��6�a�,N��5f�� ��t��J�Zy�N�a�f�=C�u�����y����b��و�3�u�6��&�郡ݕ�;���>�2C��us�s�1f7;q����F��J��ju��K���C�����I=��Z"{�x�I�u��{�Axȱ9�A�r��&Ш��Ls�X�[5��%5!#:�ߵ�'�7����e8�K����6�fU5�>�uy�ϻ���e�\��[�Q��[�������$˓�#�5����6,�Q�q�]EbPz�Sp8=�xC������Z��)q���QJC� 2F�z����߶1����b�`I=���n�����������v0������ye�sCER`���ø�6��Y,)�_iH`+Y��,��0.F��]�/�uˎ�~�ͳ��T>|i5l��ߞ��<���([����>�n}�5b��[��~Uo24l�qJP�F�Q�̠��ȭY$��κ�,�4nD�[�*l����֭ΊX=�;]��D��;٢�Q&W"���W{�qp���m��M,�]`� ��,��M�	ǓW���O����[��*��˯ouZ������+r)ۏ�j�.�l��;��Eͼ�h���ˍ�h���#�=��MN5~�χV֣�Qӱ%��[��غ����$3aN�6��T]�[;k5�(��������O�'�_�q�c��Z���x|�<�S�g.�j`*�@�^ r�I�ٿ�1��8j�R�E��)
�V�e̪R�%qyy=�n�*��=�Wդ�W�|-BLV� h���l'�{����.J�\Vܕ ��S����H�&�޿��Ϣ��m)�'�P����m)c���;5�fGL�t��}�I���;�o0j&���C�Jg�� m����z��N��a����t�3>2�����9��=��^i&�_g��LGd��Wڣ������N�>�5_��C�.�)/�D7woĶ�gI��S��<��@-��{��<f�B�f�.���{q�Z�۬�G�Y3X>��1��I�����2��̝F�8[��O\������p�<LF�r�o��%�.A�]����7b�j��b�w�@��A���zZs}��ִ�?�t�����V�����O4��_�E���c�pWyR�M�Y�<%jca��/W�KS�"m{F���+��I���ʆ�ɱʆ��p�����?��dc+'�s#�M7ƚ��f������K%�H�$&�����q��b��kz�����AXV�87Xn�OZ���wJJk������St�7�����Um�B�)����rVL���j�\lǆ����g��>(^�N910���^�>�ɻU6惽�Yװ)��| �9����,r��Q�$&���lP�\|IS��E��W�����?�����@��@c�n[�R=��05��$�>���K�1���{�[���K�CS�^��\>��Y�Q�ѿ|�[i%�※��
=��|�A�Y�=�yK��G@��0��|F�c���$nK	endh��R���1�쌥�!y�'��c�4�t?��+V��\�9p�9�)c�����>&��y5ʮ�;�8��