�4,��/���qQӦu��~���/��&����2P[�]Y(�V�RK������1�V��ᎌ��脈|-�)��^=��F����H��h�l��4���<J�1�L%%³ zu��W]��1�T,��-�*�20���4�R��* �f���G�f�v~����Q������+0æL���	��L���������y�^k��PwX4a��r=D���1�F �@����Gǅ�~�u|�r���,�(���6�c25�yT�1�`�,��:Zb��t��9䏸���B�����[�E��C�����<Z7_�)��;�#2�:��C����`��{^��ZHTd�l��q_�-���ۅ���f/P��=� �<��['=$�a��L��Z�VNn���W���
R i~������#Gx� �~^�p;�M��|���:ٲ���R!����.n������Ns[���K�Gm̅g����u&�X7��W�Z� ]����w!{�f��	�u68.�b#�XO�����&�>�$��]�ZҚ��O��nW)q׍�[$���:a���k��k�|�0�'�q��K`�y�D�P�(�;ف��rЮ(�%�a�X~EQ�e��u�8GgJ���_;ށI!�*n�h�"B�P�r溧ou������:�"lnp'�0Kx�g��ׁ&�+ n6��t��A�)z�#s�J�]N�j�?�k��)	�*�[J����v���4n{Ld�*L���k��#���Wփ��9��0=�:F���p���7{D�}���~��<ߤ�+S��F�é���Zy����	�L3M	$k�b��_�7���0<��dbo�u��)�72xl�
���v��`�/ǉ}Q��]�a�� ^��Jq�gU�U�:��N
���|����/�ls�.��Da�%k�A� �B��s�O0������-��ہ��7�gC��N^��R���C0ך�����j���sۗ�̕ظ2�ɼ���Rw��S��&�U;!�w�T��_��d����6���lD��0(J�d�I��	4�b���s<�OҦ��(���,�?�� 9%2�5�H*#�$�������0	�/��hI�Pգ�i�u>4�6��GS7�/�Ulsڷ*�3�����^�[��W��g5��g��m���m0��V���x^�go��o��Sx3,��x�gY�Vmo}��?�O>�nZ6��]5��2p��-���w|���?G�P��w�?�8w���2Io��#$��������k/WD��'g��Pկ8����9o�j����	g�lp�HQ�1u 4��Y�cۺ=���B�<MN��i�����x�t��s�g̠n�]�f׹�@�l^��߶O���ð9��wzM�����87z�y-�Mܰk�u@>7u���{}Z��%��~�3� ��3�(H�qR���m�^2���m�;��T��X�4��4���O�jO� {g��"6N�u̺-GG����O1P]����D4%
$fX=D�sV��������,R��^��m���mJk~�d�`ҁ�0���r�mB0�^�Q�֩
�p￲>@�;�l٠c<�J�PӜ=������I�h�\�gAG��ғ�`&����~��&:b�'*&��3���*����e? ox�&��k�ȏTj�r��"���l�!^�+����g�uY���m[SMm����rW�����������֋�B[���b�, G�C�aoC��N/K^8]��E� ��ꄈe\ji��M&�������8Au�^�}����!�
E��2��w�tg*�g����������{/�j����Kܦ��M������!>.Q��&»��RbM6n!�l�B��rQz�f�sq􁏣���� �9����eE���n�Sw2�������%�=�*��3N��G�2U�?��<)>L���M������k�[�d��.9@{���0\������,&�I���\�`�mNT>�F*\�<�i+���x�o�Vyi �c�}�S�e�� �/(�N������g$)���/���c���v,&����Ȏ���)�3��/b�T�PJ3}[i+}�9��r+��?JfBM����Mr�+o�������z�� ����ډG�������A�����v骋�=�݂l��Ɔ�ь�}�eyy$��9Vl�%��eA�D�8$����9m��#��s�H�T���G���j���!w��l���y���c�:��
����d.JcdjM/����M9�/�,���z'!�	8Q|߲W�?�xз1��ࢠ���@&R�)?y �%�|{؞�u?��2��k#�<'~?A�;�}n*8���_�>��k\�Go�����Ao��B��:a�T�[�(?q[��tG�Z\����y�f�đU�^X��,eV� `#VX�$�i#��l���Ѽ�W[�>h�vP����C1%.�Y:�r�З��0��y�)�B=�N�[ml`ց�Ķ�sɓ�C9�z>����4�I�Ci�QvĬ_/1L���Ц�6f�ͮ��ux��wzk�dI�L��;F �� P��Э�5yxT�h8KƏ�<l��%b`�hIL�{��S V�:�!�}������B{��&7�� ����@Sɰ?��3��+��y���_
1�4�!��:����CCs�+<U��D3�~�ϔ8����P�1�gd���\�����p���T M�@��̨C����h���<������e��e?J�b�G<�g��DސDo�I��4��]��?�mG��<9����?!�z[b8n_�^�:SH��[	�s�{��N0�+y��7�/�`�C���4~*�� �}��!/;���i����w)�t	ߍ�,�"p����^t��#G�z����Z��C �!�C!<������;�HjPbj>��b�s�5(��;�j��m����ІX&�g=�]�e
�ޅ���������^��p�߶����l�Uע�Ȣ)�ZgC� �}p��bK�hdj}��H`��~��E���qW��s��������{���)��\4O��n��
I;��7��͕��Lć�`�5�����6��U͓����v�$�B�"?�\e�2��\�A[�صoM���|/F�ŋ�������ǯ�h�▤(�����?�����#��^Q�|��@���3i�EF�q���N�D�n�#GL|$� �}B,cfUF��8��+@h����Ӱ�i�I�G\C5����!i��"h=<Bx[�
���x䋜
87�:�$�tp�ƭ��v�\�=�SD%�vƙn������-*8�?�b)�(nG�Qc)����r�'j��Dc��s����t��w��Gd5���³�D'��4�h�b�n�/ ��`F��{��^��y��y�[�W� ;�zGCϑzd���(�������L6�{����qz?�O�=����l*tGǾӁ��k(T��QzK䍺�hV�_yK��UC/Օ���:��<��O?�|=�� L�Ew\ L�܆w�`��ꆆ�"v��}:�W+� �+TE�l��I9����
��v%�2�u_NaA�ˡK�����e�iߠ8���)ms*Q���w�^cԗ,�(�@~sz��t.����l7O�h-b�f��4wi�7���૧�����R�I"n�q`g�tЅ��;i7k��xe��,��q��)�W���>܄a�&씾땗"�<7���rXNY�J�t��'ԹR�g*��I^�����i�ϩ��9�jH���{���G�P�hH���d:G�Z�0�B��Kxtg����=��݋fe��aE��OǊ"'ew�p��&�.�EuX@\J���[!x`0gw=���w\P�LٹT�@-#�×�{`���~8��U�2�c\a����Æ|��	���&�Y}S�=�BM���xop����ZK�ڜ�����DV���+{�s%C<?��� &��n�U?J�����*���,���'֞Z,�sN8@ܱ>��B��יH(֐br�7����7ց����	�+y��F���P�y��I@ǜ�C0�`Yap*�y�>B�l	3T�����̝�	���Q<�a6��9�Gc!2��2|�>�CNkҴ�ic��u4ZP��E��.o k�O�+n�ph8�(V��f���A�8�hn��JRʉ|)�=����f�K�	�����R%^���J
GB����-���M~Qτ(����l���C�?d��P���t�J^��(��\Uvj���oh���EI���}+�_'|r7C��Rxj��e����
���Й����N"��H �����ڋ�M���8����6!���!��~Y^tF��_��9�d�':衯��)�P�10��Z�
�����-�V����wR��k�D�)s"*y�:�_�!��g� �2��%AY86���YJQV����)�`p(�$E�{�Y�TS�|Q��^�D��ĵ���k"�~��3���_�ӭja�=�k��X=��9PDb��+Wc���o�a��&H��\R��R��`�6�Ȯ��z-$���!\���1�A�u�Rmv�w*-�i%�≎"ݠ�����5�`MbOxm�Խ]�|�1�L���.��`�M%��'93.f!�ιq�*Ъ�{`�P���y��W�0O�(�����ʄGf7͉_�8#�kl�U�gl�wY|+��Ѕ�T�i	�C7Z��dm�����
#)}��2C́��/��X�0%�N�d�ޡ�֖]L=�x'�0{{���0�~���ܼ�G�j��{_Iv��G}��Q�08�������v��5I-|fԴ���@��;��jg���&��
�g	Sî����b���E�|s�!��{�������z"���p0�ɿV��W�\�BaC�h����48\ۭ5��L ,��+'�)c��#w��#�ܘ"�d١L(	�Dnz �:�;���g��[�<Jˁ�����5w��>��!�E0(�M�q������{q ϲ����^IJ�3Q�C��[oxLr�^+�	o0��?ӌ��ߩ8�
燤(�#��%r��
B�E	6�b;�����:��>avX�U�©�eD�{�jX���G2�sJW�b>��n<�IH~J:�J�u���UT\��� ��C���и[pw�.��qw�q�ƒ��xC���}��8g�{=ժ�֘sT�)�?�o
tm�TE��T�/�[)j������j�`[e��f����[����=����x�í1R��)O���i�Mn[N��)O�D�I��u�G�*[���~7�5ki���jv�l��Ja�.p�B��r~�����f~��Q�:��Y{���fK6��_��9����j��m.��G���A���h58�s�I�qK�{�?sV��|$��w����� ˍCg��2�ۊ�������Jο[�#��=���`<\�����F�d���9�jX��BkT
�;�FsZ��"N�e�5|��q���e�HJ��J�J@
�*�'�G�(��AM��>yc^r(c�̲_�^j��,�w����C96 ��
�36��}ǖ02glPA�ânY�\���k�jrOE�2{��C-���HC�]��y�3�q!SF�#��p�lʭ�G�sT7�����$V𙈄� �(��.HwɎ;�����V�����S~�)��7��z��^�����Z��>Ì��'����ONN�����t��:�-륿�����H��p��v�XL����ڭ���y�.	�;g �ھ_?�V�@P��M��{<�@f�O?����b�K�2��d��bn������9!�9}�}�{��ح�C��ՙʧ�7ȕ��ݡpX�?���OՈ�Z�ҚL��
h�d�E�+�ڂ-)aE���2UJA�L[�~&MP��qu+N%F
��:���.
j^zu�j���!�Y�cu�.�wʎ��u�U���8''6^G��s\���]2����җe���O0R��Q��kvf�}�v�q�ЫEg�|��y�u�����<�aBp�-�����L�b�0E?J�Đv0I����:�Z�4���/�8����e��7D�l�]�C�φ�n�CL�j4l������l���T|Z��B�	��8�'�ӉQ)_e�P|���E�R-�G��3'C0����I���8	[E���kùϞ��²l�rZʏ6�Ŀ�_�x���ѯ��cMеn���t)�=�n��7�c�KΩ��إ�F6�zɏ����c�ۺ��޶���޵Aw�ީ�N��-�2DG�$��aB�J���53!�@��u4��hz39�򜯔��G"����K��5։�~��I5��OS�8_�o����i�sT�@-O�:�D�C8�TNRE������^�1ͽӢ���'R!������^�%�c�L�8�=��+ݘ<)tn����8+��fE��i�
D���L��h�	'J��j�b�Z]��p�d�pհ��K�t��[9��7�;%�lQa$�������w���;��azy��O�u��
 �Ё�W���|f�ܖ�S�ӗs��/��oY�
]��n:ގ��*_��N�]k���喞&E"2�6����_��"36���/�[gq�|V�r%��7�����T�ސ9����k
�����	uI��6w��Q�T�n��m��R�=�=���ux
�#\�S)Z��WI��Ak\�I�v�v��Fl\�Y��pl������|`�D�$�_�y��ԕ�]�j�)�mǊ��:��9&��3�E5���n�@�����z	�&��[�'�nx�G*[q��X8�):�fZ���'ج��&g��ȻCYK����/���Ν��),T�m6��]έ���z�6t�&q�C3�Ia����Ϲ��AW�������H�e��Դ���g��K#370IM�լ(�����b�:�x��1�ү��B�,���i'}`�z�.�L7�N՟���lB�'m��;dfO�o����~� +�36-6�`6�m���X�I4�z��vJ�Kr�������tK���՝u߾Z���g �Gg�gT���E9�3�|+�M�M}��~�cY�mp;��XI�I�B�MƍꁰU�0�j_F[[�������"HU[�����=�m�}�Q�A�jc��>�/�/YHVt�OUTG �.*ȡ$�]P_X\Xu�b����{+@B���/^��C�[���}�X FK���E#�S��*w�����*&D�֝��n�Q�:�}�i}������DC��f�*�y��h4��j�����֫�U�Mc��@���{��k�ꃔ�t�ս��m��x��jWH@b��+�����ܾ���<i=�2AK6���
bU���OA��>C� א��IH5��%c-�	8��тX
j�[�
 �]��{E'8��Be��#��y������_fN����Ŝ$k�ko���/@WEբ�D��]��PF��ȶX/v�����'de��^Ѓ��amݚ��'=�f�T�:P>�v�T9&3e�"m�<8`�zZ���_J��|�;/�����NY������|S*� ��_�\Kj�X�o?�c\�?]�k��(��
O8��I��W�ό�D�v��{鼁6J�;\ݙ�ʇ�O���� �;�uv}�F�I����/ H��i;/��U���i
ScB���ح�d�l��#�}!�C�V���R��x1�T-��k�<����ր�~6Y���x��y�ʟ���O����.n��*�f��g ���7��S��v��wK@�ܯ�(-��g�m�?x.U�{!��iB-X��S���j�L�-i��N��R�k���4u�n�
&ʛ��N��^�z��#�ğ?>���>�0��%9�.*�6I�}����'L�ղ�ƭ7>y&�M��sd��:L�lG�މ��)�m�����w.0k9f]%8��Q�qu���FD�Vՠ
nmMj��H'�ƚ�xvh=2�O&�]g�N�cU��-$����	�oȭNమ^��51'b�_B���t^�{(E�_W�c!g��9��E&it���v؁U�开G ����뉥x�vOŘ�2_��WJ֐?���؞���-0Di��×k?�����؟��n-dt�sߘ��[�vKXES4��z���;����V4ik��/�)V���jZ�P��V���eL�}���ͅ�1�������V[�\����a`�;��F���L�\U'��k�{�a���'Ι�����g�S�[�[�{
aZ,Mz�^s�r��5B��)��i) ���Z�o˅������P9�vj����ᩔsB|2�����0
�z!��	�[��+�]$�����\���C#��"ұ�D�*���w~�Y'Q���T,�~E�9p���>pib����.r��ێo�ߨs�h��w��P|1��:�5�]��[�-�M7���g��$��>Z��ʲ�T��7*=	_��FU+����W;,������
��g�a�0٨o=��?`p��0T.��X7�óݯ�>�,�	[�E��a�wLM�F�pk��������� � �n_U�e?˩��B˓�ٚZb�`��Ƌ��S��[��]-��{�xgX��T�$����	����U����U���I6��-�-�-�W}��S��s�XT2�E2����mkeOo���s4�9�.�F:!֑�w3F��g��;�=�9�<f�G��qfg����xM�G|�>�>�6V��ϟ�� Cڳ8�?�|F�����p����4�o�iB��n���j5W�:�����]��í��["�n��T���a���lWn�����C��~ ���&��R��m<>�`L��"��+!UZd�6�|�t��T�X"�e%�Uv�MXu��5Llmھ��������o[��y_ ~}�7d���l��R9�O���'���aŖLS)O��3���Ɔc����sɧT�G�]ӻ��~n�N�H�3y9[�B�϶=��
檸-��`qV�!��̠P�1�w:23�#�4ʪ�c�HԾ��Pm�T÷kPƦ��Wok|���f���-�E&#��DD��iz�z�{Xz�t�t�让hx�WGjhѨkj�2,�8Gչ�2�2F�9g�A���
��3��r5����5�u�Y�C�LnKnN����O�q�_�uB{���m�y�u��(0=�����my�̮�C!�t��c��w���e.I^0��v��G�V�%1ׁӁ���`��q�V�b1[����pH�G4K�e��#��=��ة�P}h��2� ���� =�z�a�ڑ�J,��=yf|���1������;ܫ]|�2��Y��ګU����!��}�����e�ijSv�%��l*�0Q��%2C�ؖLO�av�ګ<p^��
W�8+���C�jј��Żq٦O*y�66�D�uZ<�%X(
��ɒX�5�a�XO���Y"��3~K��=\�ml� Y�������￺�pQS[ٿ�)�mR��'ɂ����u��l��Y�:�)���9n�9��
�)2�&�����"��_�5)|ϗ�_�ȯ
����T���¾��#=�wX����7P������X��4 �O�f��$��l� g�٨�3������\ț~�t�e�lZ�4�vԭO}Pi����y�0� �CA���O$���J�a�mF�����$�c��C�wJn&�AjSM����xT�pi��+4��@�K�z��/���C�Y)LՕ�,��!��rQ���m��ԲpnVR�TKNVN]�z/J����7��f-�]��'����B���d�4Q�=))|�O��D��	���p�_�o�g���龁�Z!n��,����g�G�a��'�C�\E��\��	Ebne��h�p�0�=��q��97��̴�r��UҽG�CP�v�	�za*Z�OW��0��7$cA�)�F|U)����v�dڍ��^N&��&:Ë���R��}�d%�����eA�(��?%|x�YK���߹[~ Jf��/	����.k�EV����9Q"I�����_�B��#�q���C�sU4�Uk�]����V�_%��4Fվ��3�b�b� �D���MH�#O�<�i�j��5�{`��I�;�Ct/�h/�A���e�Dv 2�¦��h��Ū�,�H�
"���4���[������IQ3ٍ<>kn�f�~J�D�/Fl��?���~�ew�Y�FHp�M����ٔ�l��u�&Lz�Q�����_�wq�}�eS��Y ̀~��55[����];Zz�`i	ɠS���#$z]�0����h�(*+��$�3���{�qB�@ ��R�F��A^��`�*̀��d���ߠ��YVhZ��gEˣ)0I�A�V׷5����W�Ω���C���j�����3`٩���蠏�`��l�N��~��}�`��a�U�Z����n��F4�^�E?����p�5��:B
�#��2^�޶
b4r"�.S����*Vk�E�< ۙ�C�XK�*�ﺟ��b(���q�!x�>��5�V�O����:���/�<�8B;�n#��)�oOo{ ľ��12�a�yYy ��L�.���l��b:����r����(Y���+(!8��T���cӒ��"��g�9q�����׳w�6As���Pe���֪"W0�3;Ǯ�
kk�"ݞqnx�y����4;��m�+s��5��l��J�zQ��ꙡc�ݲ�F����ѻ��i�z޲�%��$�����o�=�t��z�U/j�!�,�tN{Dm5��%���/�p�� �mC/nr���l���
c��	?|���"q�_b�? ��9[Z��
�i�F2x��G[�$��cG�y��̛Jb����Sy~�I�*Dolw&m�݋ym���RSW�G��fS/�װ�5OQhRSk�ÊEDD�Ļ�:߆�_�G��\z_�zgg��A
��9!�z�Br"�г��\D�gY�^a����s4Z�/v��
U���U�+���c�n�m��K�c�L�<"V3[LPZ��M��� Ãa���-��Qb���SBH��/$�Yr:�V��:���#4Z���}�Ik��/I��VO��Ǭ���y�5���HZ�7pp��{��C�ë3,���U��珻�ۘ��h�K�3��,u��,��EJk��	��&id	�b�\�b',!��8I�=�������Љ/�x�B$�bE���~1�tl�qh�W�L>�Z�X�Z�UE�~�J�k�Z����4(�䢔��B����m9'u7_d���*�����J�i
�؛���	<�v��� P�� �e�1�R/M�cѸ��N�|��2��5�td{H����`u���z*jO1G���̃iD��G���rW�!��b���
y0m�9���PcH�s"{w���P�Rd7��V�����ΰ���*׶8|�����/!��ן ä>i��|H��4���F��G���F��a��!j�Ċ���-�z>�.&x�n+�ϣ8�C=�����)��(~}RV˰�+��H@��SSBUI�����b,�܉�J�k�$.�a�*^.q
�П�*����z��-�>�>����`}�^��ۙ6�p9����3Y*2y�31��%>������V3 ���"8��B�D�#�[���?ŷ��� ��G�����(`�*�Ch����`�N��N�a�o�^����ݘ��{�N[��sMb~\6?|A��)s���uF��x+������S�¶Xx0�E�,����_IU���ឋc/̼���/�zB�X�:j�D�zx��)����g�"`E�HG��.��R���p���&��B��˝��9�]��N�?|Ck�~o�%v`����k�博����C����k��_"l�YR0#���,��W��Cˈgry����=7�3���,ө��x��?Y��Z3Z����9�Z׸��	���=9;�<�w����&px�1H���ī��h�1
�s\�5�9Z3�f�Ҙ�>�K�9a�z�(4k����ك�uBb6H��������Gz����rJ���9ȧ�t�N;��
b���Q�
to��'cPƒ�h�y&y��:Z�NmX��!������Ne�pD�K]<����"ǧ�.VɊ�A��Ӏ	#��_2ӣ���A13�ɚ��wSQ�=�rg�u��c��.C�x5�u���nxw9HJ��	�#�#%���XƓȇ��yn@I��=#��vp��F�5g6����"f�H�v�n*���ϕ���@B{^�,���76[~ά�c<��y�uu��bYE�N����vrg��?Sw�&���9�ϥ#�ċI��8��O�1�D�&H�g�s,�V�k��d���nf�A\?V�t$�L)�Я��e����l��{J�ȼ���r����!�D�$��KD4/3�.�W�,�G}���6��'o6Q�D�M=�h��+B�=l��SP�l�#�=|�O"֬9}�*�y��!ii���M��ҐD;�,y��<�@��b��HܔY�����j^k��VƐf/`y�����e��>�Ϲ��!��'�|$h�<��p_٠�F���9' 0
љp�M��s=�U<��胾�7�|�¸��ܓ0�pݪq2_}"��)�1�=��h�쯌�B(VǖF?;���0�<3c��S�O�,�٥�1)�S�a�Y��Jp8�߭�KZ��œ�`�X"�Ґ�6^�7�3�Z�������!!0^Z�J ��W���ͼ�=��f0H:B���Z��8-�n+C�	�`^ʕĩ��b�,,�R����(�
@7r��=�aRv��8{�^��ʤ �c%��g���y�Qcu�C1�|��8�]�!�c@m�ҝ�Jb��yQ9l�/�ʠ#�/lc���rKI��r�������fwU��ڊJ���r�7��8�ʙu���[l#�"�,�O5���-[dk�c �<����n����ܟ/2�c8���?�	G�7{�D��f�#N���JÁ��o�l��1jn�E���G��J%�C�آ��0;�ߦC��@��2R�5a�B����n�$0.��@�p�Y���Ls�£G{���gB�<����͛_�h�v0a}ʐ��v�X���g����`�
��-�QH���z���2�V�p�^d~H��QN/��ޣ�T/ǳiR��k������J�^i�����
%�}��#�8�UB�8kK����S��7�Gv��Mph[�}G7D���~2A����`��)e��0�&2�J��K�4�W.�St���#FJǯ����h���)e�D9?����\�f���?7WN�*3y�������^��a=� ��w]q�v��V��p丗 P��k��Q�{���F�aR�$��J1���E��)�Di?!;	���Fv�Q��T*]7��@����ۺlkKLVZ��n�,(�����Y����r�!O@k��e7b��s�kz
ϕN���F@���K�R�O~M�F��5��Ćq����;ꎪOix�rL�1����X��1Tc��i�T˵�jd��~]����\j��k-�q|Q#�ݪ &�syv֫y�p��~�
�?���=����ƻ���O��Qrg��=�<��Nz6>�����[Cps��W>�4�z�Q�����hމy�g_n꬙��ҏ������z��Ja i�b懟��G;6��8ڃ�;����5�P\�8��@�ϖ�k�BSM|�XR-A�:��+�J���
sP~�cBV�Q��9�q���7���eߛZ��2�
Q:�2�~�d����|��&�Ao�F�����~
�Ȃ���>�W����v]�+�)��|�ǟ'�L��E��[=z���bj�h:����Q�Q�u88�_��샒��^D'Ѿ�P��m���܂�����U�Ơ������~���?���ߪ_~�\-���M�nw4"���v����)��'�/��M�aJW��e�����.J07���&~dМ=����JG��OAw�m���~��+H�K&[j4j����7���u*���g	��n}g��8?�G��q;1��	��}���Cߜ鬻���i�}Oޚ$�,М�%��������oaA�3�j��ӏY���������CX��t���?i-2�H�3%G,YNڙ���|����k�Lx�b���AՏ��!!��ť���>������^W1�_��ǂ����X3O���*���7B*!U�a-�Ü㫈�6���E��y �