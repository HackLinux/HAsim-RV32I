������ll����++��������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������WW��������  ��������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������bb��bb��ll����������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��������������  ��  ������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ������  ��  ��  ��  ��������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ������  ��  ��  ��  ��������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ��  ��  ��  ��  ��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ��  ��  ������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ����������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������  ��  ��  ��  ��  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������  ��  ��  ��  ��  ��  ��  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������  ��  ��  ��  ��  ��  ��  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������  ��  ��  ��  ������  ��  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������  ��  ��  ��  ������  ��  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������  ��  ��������������  ��  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������ll��bb��bb����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������  ��������WW��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������++����ll����������44����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������,,��44������������������  ��QQ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������������������������..����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������������������  ��88����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������II��==��������������]]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������''������..������//��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������11����������WW������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������WW��  ��vv������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������xx��  ��SS������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������  ������������,,����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������$$����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ����    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ���    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ��� ���    �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���� ��� ��� ��� ��� ���    �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ���� ��� ��� ���         TRUEVISION-XFILE.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                < K  ��� ��� ��� ���    �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ���� ��� ��� ��� ��� ���    �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���� ��� ���    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ���    �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������<<������WW��������������   ����    �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������((����##��������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������FF��  ��QQ����������kk��  ��xx����������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������__��<<��������������������<<����������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@@������&&��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ii��  ��FF����������``��((��''����������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������88��  ������������������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������..��������������������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������MM��  ��xx����������������BB����������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������))����������<<��  ��{{����������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������CC��  ��������22��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������{{��ff��bb����������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��������������  ��  ��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ������  ��  ��  ��  ����������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ������  ��  ��  ��  ����������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ��  ��  ��  ��  ����������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ��  ��  ��������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ��  ��  ������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  ��  ����������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������  ��  ��  ��  ��  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������  ��  ��  ��  ��  ��  ��  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������  ��  ��  ��  ��  ��  ��  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������  ��  ��  ��  ������  ��  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������  ��  ��  ��  ������  ��  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������  ��  ��������������  ��  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������bb��ff��{{������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������22��������  ��CC��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������{{��  ��<<����������))����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������BB����������������xx��  ��MM����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������..����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������������������  ��88����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������''��((��``����������FF��  ��ii����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������&&������@@������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������<<��������������������<<��__����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������xx��  ��kk����������QQ��  ��FF����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������##����((��������������������������