�g!@�`�p��9qf�A����6��ݜv���G�n���V@���}�<�5{�u�i��b��	Q�1x�5�<Ud@|5�ҝ�į.�=yX<�+�WOπ�9j��s�#Ө���
�)�.��O:���oTEMP������F�eG�n��G��}� � R���5�����ő�e�F>��W���#�26Nx���cI�=/�q3�`y!�����=`y�/)�ww�\.�at�^��S����H�sX����TA���aL�َ�@Tm��Tt����V��f6�F-aV�~O�=4O���˶��(�p��Xf�p1SC������{tЀ WE��m1%Y
�{Ԑ�F�V�Z�E�=���Y+�-jr��^�ekg��`�B�\F3y%N�u �O�ȉֹ��];�<���j:�"�!�mhhI� �� q��C�5v�MG=z�>��1�V��[��~��� "h�Ψ���n�Ɗ��h$�.�g���mIW*��Ǧ��� z���D�冷z$����t{a��?(�9-�����@�j}Uʏ�UF��˫�����89�����x��N��Oc��v�wUP��lT"�0���w��cnw�9�@c�PEmMF��0md&���21M��1b����P��U����H�&�`6`ڈ����0+1��T��������z��I8���"�wSe�[w��R���p��h�P'�Va]"��{��ψ����q/LIE�ҩonh5��[���NL�q���<7�=����By}�?*7�Q�b��(�so��7�����XR���f�����	2�D�����X���&bq�{v��/��
��Ã��`���G�{�J�&|��3|��Ъ���&�u:��Wa���!*|",\��E��j�����J���]����L���u�9Z>�FN+��L3..�
SE,�M�}I�ЏhպKU��SVc~F�C��_�B?p!��&f13b7mK��Nf�e�ʫ��C��G��Ey����9# ��	�~�ub��_���I�E��
Ɉ@-k<��_n�&�����&:�bJwO�JԷ��U��CPD��OX Q�TX��B�@2)�����!=�9�<�͡ڷ���Ok�$�:n� r9\> "{j�x����P��"?; E�����I��������������\�?�ņ,��6�.? H�����N?]�f`��E���>���r��Fc�\���r��
3,��0��ˋ�'�H��>G]����0[�_�K*0�G �p�GZ�}ip�"�V�J���|�s���s�p ��~C-ۺG�JU���׉���Nl����Xty�����A~��8�A?���200��驪���� /Y?��q�=������)**�	�#///%%���IKK������GxVPP �j����������
�[rn���/^�������`cc�����cgg����h|||<<<���TTT�4999�X~ ��YDD���+�РH!!!-uC++�Ș���Ư�3
3S�S�󼜃b�2#����Gd�'���tK	p�&;��z;��l`�u��6���K|���W� 	X}111`�^�|	l`���(���2i�����,��?�K�Z�����毫�YXX���R�+�t���<3���?7�����j>޿��y��rY�W?�egi�ly�X�����������ᖝ������w��[J�]\�V�����4�Y����/�����4����g�v�7�U�-fx�����p����%�q���}}�l�_Q�yg��%zzz`G����״����^��O�HCCӔ��X�RU��U��x��q\7�����Ժ�{\��%+�ꍓ��K��G,�����d�dZZ�dX��"��KEE��5��5�����ϝ��c�ݝ�ݝ���c���)�;-�'$$�(���$�x*J{J��  `�?��x��#������z�q�P�n�x�	�*Ǜ���/��:	_2&�KK���j�L�7��k&J����-:���>�[���T��q,��jR.����`���ᡊ�h��<�,H;8&����rI
q�������;_	ϖ��B���g�Ep-	%��Ҡ��⚿�5]�
H�l!�w�#�Γ��=���7MS=���W�=f��%�#Rmu5x����0!���f���*[�����A��#C�P��Y����������>���۰�룋i�� ;�Cd0�9-�2� O ���?ʞ�L#����ij�[���\x��:0�nf��P|�={]���z�jcc���y�����41We������9���=����P��&@K~l���C �;��*�@|9�[��K���-�&�OK-��!���9�^�_E���]�u�a�:��@sk����׹��,˵�{~K���[D>91�^��݇�)yR4���s� S�Ꮣ��7e��tL)�=�jWH�_��9�����H�Ðd;�o�C:rV��3z;%:b8���:ޏ�vYp�t�A~>�"[�����ɞ-:"�����1E�Y�ym���uz~��r���V�$R�3�<��^=gL�mz���T=Y���rM�����;,��r
��N��{x�35���7��/Xn�QTK���J��N�'c�V�o�&�_xGữwIĵ�r�lĵz��*ɥ��}:��l���{�o�:�HP�s�{�j�rv�}�r�yp��w۷zp�.�(���M����M��?��U����cy��6"ح[9?+z{�W;�6�Gx=@�_wR�x`��m�|�rC�mP�Jiڻ*ǭhթ�"�M��nMh+f���r���ƴ�{#��9���@�=������?ҟ�L	N~G��t@��z��eS�D�-+��&= :�J{Af-!�U��~�v������Az] u���@ɧA,�W����Ϟ_8���Ca�|#>��L��J��|�g w�Yd�����y��`Ox:9"���=	�x@3A�B�&_O�в�׶)�Yꩠ���S90�5��~(�6`TE�U@�ώv�6�Ez���ݾ�"���|ZP��q<��$^�QzN�x��2S������K��y�5H�p'�c��� �ˉ����e$�[�q��?�H>j�Dݩ�%1��}�"q\P灂��[X8^V��}�٫E��;��XW-�ktZ;rr���?�w�������0���\F������7���պ�b��~%���F�����Ѡ�����_Ժ���Z��7`ہJ [�À��� w�P���Y�ar���$5�v;���W��_L�-��2��u~b#1�~S�G�꧂�s\�N����T"�C�_,��=�{��]^�=[V���#N	��N���Z�;a�����=5Ԙ;X ���).�J����kV�5���D�!�X|	#L�H}l�� G�m�)�f{���q��W\����T�20ѻ�̅g��;@���T�
���<��^���o�jH������������И�?�M�V�����c�E�K����ݙ�a`�C=n�K�C�Z%�tY��Y�*	��F��g�>'W�#��{�-�<]7!E�|ׅ|G-L��s��J ��CM{�{���N��ꭂ¼k��.���[�� �H;����:�,��,h��bF�~�"��p�N�?�ټD)�M�n5_�h�\��'�pm��6}��6���3�ԕ3�H����ֲǕ�z!u�j)�����mGgN��_h�T�4څՉ�� ��]W�˰~��)�OJY7��.������YY�I�OP�.�A�aQr���j3�	�4��˦�������_13�<�૟�#�~_���f`Iv��R���E8#�}���ző8'���e�`Ш*����I�V.�������k��3";������I��k����{y������ɢ�7gR��y�}we���'fs�(�,���Rn>����sxȸ9U�\ګӛ<�m�,ﭒ�[p��H3YPP0�|��@�Kߒ���{h�Q�/�[�����:�Nu�i��g�Z}ƇbC�w��tџ���j���Q�dz�7�Y��3�5o�F���ge��P�����.�	@���S3/vCo���N{�^l�su�0o�R�W=X6��"�b,^;�{2g٪d�̂���xL�X������Y-��{-zh'�������'O���5���.�o���m�n"�`gI�9��7���2ڑL���5��|�\ ]xg�Tu�qX�̆���{y=��KAm2/�48�n.�}t��CE����#�
��,�nU@O��*�r�$��#��|�ӣ�"�!��<X����I�s�E����H+�u~�>꼸`ZV��{;���:��Q0�C��l݅�ؑe6Pȋ�ikى�E��5"���+��� %�u�ٜ=�~^��w���Z��f���͍�
�.�X<�=gϷJ�Z�>�}�vkܮ�`N�����)�������$�4�����P�~A�X&���{����;��M>�Q&���G��:�о��r��G=��k9��e,�P>t��U'~�	 �$ml��E����$�3���T+�;�@�K?U<��&���M�8���N?���k陎�Nq{Y�
��B�D����I���<�~�ߨ֬�*�b�Q6�y܍��`�N����Y����\2�	���w�M`lA����~%	�N�$4�Y��C�(���`YS��#��+<P�ϔ����� *�?�e����6{��-nAG?����`@H�姁t�&��
�H5 7�rrj���}��� X ]�&�7v�j�D�sX��ǳ�h ����6�p�?v���U�����7�����oT��\`~>��k������u]���T�Fj���S(��p9Oj�z���*�H��� yp�,����%4����?4��-�����&�>e�W4��ό�|���|!@��@�A@���ti� 0	>|/��;[��R��Mkh_M`�G���Rm��Ė7��Vt�/�-�A6*�o�u�������o\�R����. �;��OT��I����zs�T��w�%�?�QA� y�����$�7Q�.�|s�	(\�WE�i����&��J�>+����d�����4q��}��ҺK�\1��#�R�@[�|�Ą�P|cS�-[`dO�n`��g�M��jXxǕy�]ݜM+X2�J�"����͞i�s��\�=;g���\�Ȅ3u����?�Ź{s���5�\�� �+^�p��{��&��3�+viI�[�jE�A{!җ�ٸ�[S
�"��F���P KZ�r�M:��5�w�n���;ŦX�
�@k:80"��C������ϱ#6��|��0��9GN6)������5ף���_�3f��QƮY�UM��P���q�I)��É*��lt..��vp�>pi�����?����U���IH���/�*��i��OP׏$?=C��������L�>}yEZ9i�}�
GU��:|�u�3X���n��|��K�3��o�=��1��绕9�Ѯ?j�ISA�wžI�Ԧ�w�`?˰��q�v}�Q�ir X_���k�b>��>ӻ��=#�|���M�����H^
�9����۱Fަ<�p�0�� 1g��Ջ _�F
I2�s�`+ �8�iҰn!/�`V4�@q�_���E�y���a�o؟��珙��4�F�^�X����i��brt�n+�����	b�?Z5Q�|��)�mXI�#�ʂ�!��=���T���A~��A���`��/�{�� :D�����(���<l��⻥��7.p/� �ޝ���dĀ���L+�G��!�W跿��à����{��$��͹�p���O_��7�ӧ��!���O�Q�����Jq�'=����q�;�3g���o����D�m�a%���5«�ƷL�~���L�5�C#�~�o�ys�'�-���`0�#%���{������A�9�z����p�
t-	Vң`b�[��Y;�sdj�ʰ=���v��pk� �����g�Q�v>&md���.��_�7�5�h;�@\��_��@��2-r�Kl:��6��}�xG�����k8��_���CD�GJާ6t�Ho����m�V� �&�L�F���
[VsS����p
�ێ?,A��H@��ZG�q��vK��;�N��מ35� yI��Ժ����d�q#�oCk���!��Uъ�l��%�;�I'�P���;$���@�R���p��Eup=
yMe
���B�Q��m-�J?�ˊ��zθXőBrJݪ�� ���;�a<��Oa��U�.�R��� ۨe��9��$dKX��S4�eh�?9\\)u�ȸ*_`w*�I�(~QϬ.S�0T ��S�Q��@�D�4D~�ް`��W�k�������]˽<�g���\��m�&jh@7��C���G�{�>:�F�r��nkP/�1pB�/0���[�+����{���Kp�A=/�Գ7�i�=���";`di=�	� ������i�?���Y	�g�˲�<��Z���cD�"�(r;��@lj���/�j"N�77�`�������i�6+������x�d� >�r���S�����-<Ӣ��m2@9!{�",�6��|>n8��X'����BB������X�k�e���+��|��Z�S��?2v{5����V-�m�H
�t�$+�������@WgN�[2�7_����_&^N|�a;wq~(�]�H{���aǏ�]92
��������h�"��NS���8�C�&`����^Ԗ�U�=d���mc��{�)�'I�#��r���w����1��W����������������ϟ?����xxxXXX?�߿��������������~�:66VRR�?GFFNNN�֣g��S�+0 (84,.$�3xTzL14
VtJrd8lD2$�Xl�9Y��II���^�3�R�s�0		�~�?�8�Nee}�"c����~nn~~�C�	  ����3w�G��g�eЯ�a��F�y����{�`�x��Ч�VE��u�Q�7ލ��%N�3ܦ3�V��Y�o(���1��K��6+A�!�A���Ƙr�7h|�8�j%�YJk/i��X��a��M��ކ�JW�&fѤ+
y�8y�Q�Ӷ��v:dw����h��6;]vg`�����P�U�@�f�2�b�ŏ�.e�Şd��)�	�QE�����wzF�ѝ�`�|,T��
&�Y��&��cPz�Vkp���/L�Z�U�'p�<�L�u�[�^XΙ�#���90��I����0�8�v<XT��$[�1��"��I/C��\B��P�&!Z`���!�9M�y�l�55����(��9a�m4�Ձ��S�k�������n�ޘ؍3�{�Sߙj�"���̹X��q���,a��*��^����NA����6uZ�,k�>V2
&���+qDWj5�v)��S�րg�B�q�,�S<��0Vi]����3�����3j9��za�S)Ak��?w����R���;�lـ�r�
N}���y@dٚ��pjă������cDZ>��UJܳ���uc�D��;��F��|���և��ևͥ戽f�w-��K�ݘRzg;�/��/]X�S%ټ�l�8џ�wJ~_�%��g��ܛa����"�MΙaS1�� m5��I��u�����q�[�/���఩�V�Y1�����D>��.��]��u�,4��~K>]�_�3Ѣ�V��cT�뵯�D���s	u���x��RAzix���k)E�4a��_�'�|����L��P�~9Ǒ��9Bߺ����X8=v�\e¢�^E/��a5 �ɵB!0��*� gw�����L�;�{+`��<g��\�;�@�;�_On�+�Ǆq����9_)�z����t����S�j}��M�'h/M��gƮ"/�n~�`"ջ�x�8��Y�9��O	��M���������?���m
z|�����,.<���&��E�3��%�Bp�%nz�Pl���G���ikW����wz�K�2���R��VH@4q7�+��B	�1��V�����w�W�6f��U�Eh�%���Ȣ0���k�������K����+CK@~:�gt�V�G�Rg
c�߶5̆���
b��S�ߗ;$<{��{���hP.�^�������]'7w�m�vE�{l���ť���߾)��VQ-�ȋP�'HQ�IH)��e�rH$��|���h�ׯM����e�����(Է����:p2'K��
�KдAl��@�8]�<�7V�T�dLd�P*A������4g���56�
������ˁ}�GȻ��⊢mQ�`:>$,y�,	�[��[��a1Z��(�gK��	4P`*Ќ����B'���֓���S��F';����^cbb�d6���$؏E�]Q�n̺*����Fy�T�5�۝K)u��n	�����&̙#2��6;�,"y��y�!���2�]�:4CVlq�OyT+��a������a4+����ml3��R��?Fn:ԏ�j� =�V���N¥��:�y���{w��<�e��dh��\�'�"��d��/
�r�6¢�,G���ɺ���s�EH6k?v�;G8G�����1r�-=��6"�'j	�_P��k����NH���>�q�SZ�[7X���(cj��@�!0�$�f��-Ly��W����J�Riǿ�#�����o�t_�7%�~��3�2	"@LgC��30&��Z�"w�%%�Wg�CM�:��3dl�	�λ�>Uq��n�����R�gA�l݋��1��Q���X\���y�c�ߘ)9C� ǝ���%B��R>͸Y��#\ݷ���J�n���kD������%UD+�е�W�Wd�i�0u<�ikqW|������G�tث�o��v�oZx��CY�QEO��ټ���-J�(�ʟ��>�=�(!:07�Y��a!�����^��&'���:���@�̧��.�VD�Bc�']�"�0�׍�i}�F5�m�ĕ�z>+��Nבd��'1埫OͧR�9�G�jԛ>�8�q�i|#���H}��f[��1��G��1��M-����}�}�\���HD��a �P��:|]d�J�?;҃IF�D�6>����_R�] ��ëT��/�F(�u��5 ͘ �^>��6��֘q��;�~:�O����a�'����ْ�%�����x-��as���$�A�p1��UK"7��be�_+�^]���g�W���Z��[���oI\~��zdJ��p���(N��k]|�t)eޡ��P��x�=�G���޹�I ��|\6$^~|���e��pA?A������c�,��:�xO���H7�Qj������Ί�ŏW�I�IO��	"~ݣ\�b��/�T��x�q%�ī�fg��]}E��U����+((

����������������0)����a@*&&&$$$,,������o(��W=�6�s�6�H�_���\�ID�~���Lh�#-�p�l�Dݤ�X^m���t���!u\�k�Y����b��gڵAͱv��1�Gg�}E�hA��J-����WOO�����?�,y{g?��XX	C���<0��$&�}��:�DU�jr�]�D�,t@@D��eu�E�v�����=�}�D�p�X���[�J��h�|���դv(I���Z=����{�Mf&o�M�� p�����?����'u�=4�#��c���	`���������EEE����5�i�u0B��$h��-�;~rٕ2��.���f���[ey�n\�Ps8��	�mЏ�[��L�1$;H�)��ST���_t��GWK�x�1����(SS��T����TRB�j�^U(H�V����
d�	/�cT.�M	��K���lщ������ �_ ���3���0�Z��R�>k���O�߬��[�rq2�#�n���w�|�{��.:�g-��/�{�
x	U e�Q��`�$#��z<�]�6c]~+\^S�ތ��~�W�=y��H�hn��6�%��1Zu��_>6+?Q�������e�3�k��`���V��)�߳�g	�tv��;[�_=h��5�(>����
5�Go%3�a���.DZ��L��@Obq(~PI锋��A��U��2�_���M�.��Z�.�mp�j���Hj���C��}wu��p5�S����W4n�	9�e��:��l��p���W�}��ư�e�U���@}~���������ͫ�\鶟4K���������G��xۤA׎���%�"�p^���O:ֻS�Z�|�o���>}�6��L�,lM{�c�ȍ���+�k�.%?!o"���o�t=62<����*3�.�3;;�>C��G]&�/�:���������������d���^���B�Lf�� �<�%o��Y(�r�gE]H1J�`j�sC�
5����'U�a^�L��u�L���@�EliQEWF&�b�AWW���������*G'�q��ĳ�B�a��a�4%�z{� _~1!X�Zm:�<�+єM���O�7v�o�	���=�W_��nd�Vf')^����5CJv�"���8�+�Pb�I��K?�ê]}Id
r-�fO���S�"K��e��\<�wTR?k����x�#�{w������l�N�P��K_
QY�ʑ�~W��b��5�eW��Y��}�����pc{h���6��я�}�)�
f������ޜ�R6_-��zN$׎��
~B���p�+�ϳK�g���
1ڗ|/_ء/�_P�������W4x�t��%&��檕�]~��Z�Cl����7�i�8Q�	;c&b*�=���� 7{ptr�2�CF�c*;��=Z��f6=::c=�&��x��	�B~:��Zt
 �J+���bź��EKj<�	'ܖРM�'�'i�/1�˞�i
	��I?|��R��z�AY�z�N�����"�Z�ۺ�W��D�89_��<�uZ��~:�����x3e��ے�p6V�U�AkY�-tg�.܆w$L��9%�5�[hõl�㘊��7?�����7������5���(,R�_�	"5�iԈ4��r�}	�� c���r�I �;��"){9��O�o���^�L[9}cy�w���w�GK��FB����3Z�ۨ^>�	H��>�󥿥4��'B���%��S-Fg�4h�;P��|�@�Q�!c��V�RőJdh�Z �.L�����f�4x�Sps2Yc}sšg���<l�f��j1\s�ǇVl�W���ߘ�������*�����TV����s=��b@��8��8[!�����<�Ϭ�����L.K�w61q�������A�j�47�CLӆ�K�H5�qW��$#e�K�뇾�o,k��q͘)*�� _Nc�������t��C�nw�l/�T�� ^��T�H�r�G)
�-�p�`���B��{(y�+G�+����?������B@\v���`c�j��g�)b�RpO�۝p�rP�vq��mk՛�%���������ܨx�t���M4�X���;Ɍ4��O�Yt����%� P $���A� @�;^��%��X�bJ@gr�����Бֹ6���$��f+.UO[�7����W���$i�M��<��<Ѭol���⠫��	! E����R����@�GMMH��������痖���'&9j����U?�$v�.x�/�V-2���o�`,O���e��,�,Y�t�g��j�q����p�3��KC첥�g�a9H����u���q��W!-/ڱ��@;�܀����(ޖ��A�������������ݟWm��,��,�h�ax�@ZjJV��,��R�`��}��R�@Y.�W��&�h��<O�D}ʑ�=j�[��?Zز�v �A��kh4�>�O����Z�����:�N�Bp�bjt�����O,����B��/غ(����`�
9��[��:WI�`F��"��?U����xzTD9�#��*`���a��E�������r}u	ai5n�����c���z�jI��4DV����hi���Gy�Auzo��3`�C���S�r���oN&[�MgpᨙI������n�~%$���� A�|�S����
W����Ì� hp�p��1�KL�3�E3u��Z��s]w�5�W;	��F-^����&"z~�����B>
8������/�
����G��5w�g��^����x�q�������8=�(rW��)���6*x�S�z(A �2+,,q.��58r΢��V%z�E}�E�{����Y31�a����{���<l^��6�w+�P3hN�����: -�a��B>������5�W@�2������(3����<Z� >�b�L�f)�n K�1���RU��2��ի%�f��3cO�&�N,���"��� 2�RG��z��������21A���B� I��}P�8Zm�qqq��G���[[[��ш�K��ꃴ44����oo�*�����9r�Z�NJ�7o�Z��rjjkU�2վ}��Z��F"yg;��777�gjj� \� ��n'r;���~�E'���΃����P�/�kk/��b[v�,�X�������e�����V^��T��Ї�s��`���#c�A���дQ@�(��S����Z#�/���cQyi#�/^^��/.f!�ڔ�IK'AԵ�d���+��������\���k6�������g�b���m�\@����EM2T����5@Z/��BZD\��e_L�o2
$���A#�I����eR�}���y���V��De�
�� R�j�9��L)���M �0�L3�Y�(��i����6n�F�gbs�p����T���&�j��Q(��{co����<�uw||�F�m�0��2ύ��9���l�2 @Wq�Q�P�9�"o���{K�Gݖ�GGG+v��HR�\?���I��eK�yA��GY�J;SSc
EьG���+����N���	/�UG�d��(�(]IA��P��򺙳`(�ҹv��A��[@�v�0��������`��5�-���g��^+.i~dd�2�܎���������,�"I�E�2�	^��p�&WUU	��A�;��p�������ut���=��WV�>}�x܄m�c�(�G���:�pH����>������d���ܙ����*���!����&�)ۏ��YEΏ~�M�����6�fJ���k����<��F�E�o,�un�__^��fjh>4v���9�S�HY�P`�0�M�������Q���@��Y��ꛋ#�3O�Pk��:�|U�� �a�n<.m�wi�/�8�ϕ�>�$>�ݨ#���^i�:_֪/�v9o�[�.�%�^I���w����f D�Z�[�4�`	�%o$�Ƞ:a���9`�9�Ͱ����r��^��wBѓ~4+��0�`��<6��u��0��ˍJ�J�i�G�D��0�<�.��p�64�4F�G�[O�s��+�3S/{���zt�i�i������vY�'����C؆�ݎd��8�}4���2"ڞ����Y�P��G!-���c�܃�o�*Z��PPP�CHR�A
�s>�
JPZ�eua�j�����0��ˉƒ��P��0�I��Y�guǵش��h�$�X�_y�B������
����yq���H'���p�C�ˠ��m\��׿���j;d�J���Z�gf���0����`���|�S'����I��͓�m�'�siҫ���ދ�<�b�z��?�\�ݏ\y���/�(u�߱�Hv�����S�J��-\Z����I��s�s)&���=��Ǭ��'�~Ӫ~p�w�>��������a�xm�ˋcGV�X��VM±��5ӝցt2�B��{~u၌�#�{��6��Ma���p�xp�����r�����:z|EA��މ{�����q�G�	\V\���O�ƹ�nC���wp��#�#��->�T�$N�p�,��]�����x��0����:d���Q~��ۺ�yR�ԇR3onӇP#?�G�Wh�ؽ�Ee��sҵZh
hx������uH���,F����|��f8:U�SE���)"o�Y-�Q�l���o�c%_���ev�cM?)w,��~�)B���o��N����Ǭ�n�m���J��sT�������-1��݆`]�#�Yե��ˆ���w-��$��f����L�S��Ua�5lv���ov�d ���䵐Vˈ|.`F�]!�fE��a;��MsA�!Ϛ}G	GSRRv�Y��nͭ�K**��H�����[�����xF �ܱ�֛1"�b[Z�{J�b!  棭ll�!{.�VhI�.�\��IŢ�熜��|�r��DK|�zA�L8���#���ʞ���H��ّ1;��9��r؃UFscn\]��!�5�M3�V���8X'#������1���yP�k��w�u^���>��m�Z��׎�A+p��-$Ns��dE��cj�� F�ǋ���9-��Ew�2����8��������a|9����D��E��Sg��j}0���̲�~%�'��*6`s�3���=F��OEYyt�8߿���|P*��#ŠcV�?�L=ܤ�:�J�$45=c�F���.�V��~vV;	0�΍I��Qk��@	�����)��"?�%~?��pPM.�:�n�a�̤��C�A
1A�0�dc=i]W�b�c� 4��C�n.R_���7ײ����p:���t{iOEMWL�j��'�q<>,�r�z�6�O	H�N��u�C��|��B�њ	���#|��%	�3�kkk�/it�k�ai��'�����m4�H�v���"�=j��7���~�J�����j�;��pd�T��M��U	+h,�]�w�z��d��<pV-�x�/'��FJy<�Y�g�b�t�
�r���<h�U�ã��h�����ᰍ��5�-Vy�r�|F�^m��X ��V�,��F�E�����w`2V��bj{�b�LOJ6�dD���NOʐ��tnm��}lb��K��&���$��=�9s�2��b0i8�Y�,�poc�r5�[@�!��?:5�/�h���SЄ�����щ�Z/��JK�J�?�i�!9sXӚk�|<:�R�v�5�h����^eUb
±Tg��(��#q�-9�P�i��2v��P�Xr��}Lz�꾉�BO+P�S3\��nT�ht�:��]��{�o��8p��<\�RgR�m5�Q�*��q9?&)�D��bG���R���;b������_��ɳő���ٟƎ�E��~��mmc����t!A�w������T�߻A<祵�uDqw��
�
�FONM?q�NNr?�!~��2j������J��؛�O_��5��E	�͹�6�4����3�����S��.]6m���>���L�����~!}�L�YPT���v��-�d?i�HHZ��d�R|�R.&���X��.&�e�M&<��k�0n�e�f��ke�ˑ��U�S�n�4��[��N��|����g�Z�T�J������Vr��]�����PACR�	x.����z���{ӇHn���S�escA��x��z�H��Q�QN$d{?\�a2�����������@ Iw��'R��2@Fp���Ciᶕ,i��/Y�[��k_���������I��R9�b17E�	1�*����뿇�>�;���d�>�=��.!�ݟ�I'���e��]k$Lܷ���t��7�Ӵ�c�!�r�^�`9z���!�9�߈�LQTH��O���Qқ�mh�C��5�e���i��U��B�+b�J� u���ɧ�"�/QgL�Z��@;���]�ߙ�v����Sc�wY�i9�M�*��.
�Ʌ�1��6?��7�J�8iE*sB�k�������+��
u��XP>l�2��q���i �Ę��2^x��$倮LP2qx��d?e%�p@�
��W���f��kL���{]��~���KN��.�b�cg�Y}�h��_�@>�%W��w���	A�?�
���������j�� vc���o��<.Ah�W����߯:�t��9G��+^'�~���?��`Q���zy�AK^� Sf��Β��mЕ�p<!&=Dģ��b	�G
�_�*,O4���,꧄~W�?�3Ɉ DjcoF���YL�%R��d��;+qnϭ��_�I�{;Lz��7�T�Ŀ�s�e�ge�`f�?����\@��@��x½?ʪ*h�ÀO��HO��Q��j�!��V%r��{��������5��'����p�o�͈�W
D�bL4B�|��
ٷ#�H��T��Y���C�(M�_*WF
H�%����30����"9�iN�@$J�]��B*1�7:ڷɂ#Xޯ*��	[���w�1g/Y�RnU�[��ϙ��������]V��H9KR���*6ф�!3��(�4�}��Q��M�ڙ���0��WJ�>�*0
�T�>��*��ND�
h]�/�&4������}n�.�h�]qcM��:�:m��BHUM�:Ґ9�n_4���ü�}�1��d&7N8�y��TgNQ�ˆM[�V���� ����B���&4+u�"zW��� �������`P���g���^#�_$<MW���ΒAp�q]ɳ3�A���8�����<xp�.��l�2�P3���3׊$ʺ����b:�[B�r_Q%:n�Uv�	�7J�ߌ��'ǍG<G�C��Yw���a��݆�^�?��ϓ����殱~�7��ޜJ�W���9]����Cf	�nۑ}�l7o�����b�#,�9-e�";8�"O��5Ik���!<���7ޭ��ZZ��V���հp�H� j���a�Z��;x�;e��1T®�G��ö�b��?j0�m��Es(���s����@�ǘ���S�	��%�k�?y�7�Qw��M��,�ȗ��{tĳ�chjM���-��K,�.Ħt����ul�?��m��s�P��w�����V�r.Ͱ����,R8�şY~�`W
5f�_\��+�ō n���$�b�$�ς��]���gY�E��^pgl�j��j�J�R��L&$��"<���\΂���6��w�Mq��(
09({r��dv24����p����D�Rz�����|#�c�)�!����t=n	���� ���s?($'1Ȕk��d�~E�\Df���9&$mf}\1|չ�b�Fc�A�:n���XbKX˾�}ׇ�wH�S��#�ՅCć����~�n���N|����P�B(�ܒE�9>9 �v���0`eG�P@���1MFP*S�.��؈O�#XZ��%N',a���{���`˰P_
P to��R���y��o}��E5�1��O���pL{H��mY�ԡK�I�6=���=�Az
a�Ñ��]��;Q�ڲ��������-��塲&$�W��VD��|IB�\.O�	�����E�O�M�"-�E�k4�!���2\ ������E.ܽaσ �I���Bx��i`�N���`��B���;� W��,����Q�b���[V���Y�L�9�"�_��ƹ�0�<� �Q���P]�\B3�" �^�8"Bj�S�p�W�	"��g$���v�6��4m�^��m! J��ޫ�
0����0I=�}�^��΅�%P����x)��4�y���6��»�S��?Z JX�g�#��ݰ�{�U{�O���r<Ǆ�|�,#ձ����? ݈���i<N�(ĨY������R�>�NT��G�_�����٢z�+�K/��di��c����0�t��4L���XȎw��ߍ�������0	�-���_7ͳ�����[�*��𨏛�5���6��?6ͤ'wY �R�����F�G�8:�5<�YΙ`�E��C��[0P_p����YrdΩ�Rp��nr6��U֑D���.8�*�����>��������4�{��٢Uw�1���p�U p ( Z @ ��q��M�M,��C=u�Y+WU��MO� �_`��S�W�I����
U��܏�K���=� �;��G��2�	 bJ��̃X��A0���FS�҂�K�Å���!F�Z�دʥ@�.��&ٚb^T�_٦�^��s���p��o�������pD�΃/A	�6�^A�B����s��l,�Ǖ߽sN�_�A�f��r'.��i�L����JCNUmm�PƼ���)E�a%�F3�Ӑ_�#,��	u�Uu�{�D2�o
;�E2��:=?���p��	^�i����:�����~��_(���۷8��c��P��H[+���;���'>��A�E��X�E��e��	�8ߗ�5�U����O��  ������i�G�g���P����i�Ӏ��Y� 4س�u�	��D
<2m�0�D���2ΝD>���N!#Z/�͗v:#$�{{{c�?l:�0�N4i����F6Z��Q�,���*d�x�J9��{%(��v����/��?�	��0 ���>罆o�(8]���ڠ@$���-�����vi��`�*H��x-�q0�Yh x��CX�/����g�d%�$����Ϭd��m��a2�=x��
Kpn/H}�,��_U�o�b�Y's;gs�l�M�W�A�	�c�>"~A>������ھg���Pf=폘w��aqܜI�3�6�/�M�SI�� ��趬���~��K��fkk�S7���}��x�HOҏ���y��;u��.�8
X�2tߣ��_Q����Eũh�q��! �ǤB�������j#����z�
Bk��K�](>��q���Y>)5<��w�8�~p|�z���ܚ����~�6%�+��=pnn�!֫����T�r�]Oo!� �T�(�2>����N`����>�ewwW��6�&�$������.`]V����9=P����"��z:UXX �CK�X��7�Kwww����twww�4�4�tIw(-"��-�H�HH�  g}�߃����\�\��fggg�[wߟa�,B�P��A�M��-�F��r����o�p�w��fv�9��V�&�Z�s\ll���z�Ù�A��^�J{�LOO�`� ���S�oU\\��P�0�#HSSӺr������*���S���\	�"Sj�B���;�������q������DC��ȸr,,,E<�9y�n�T��j����=�&+:1u4�1	t����_�z5 y�Of��::2Obbb���ȥB���+�
����}H�#�W�]�`N҃�V�c{졮 u�|V���\�36\=DC���R���$5�'Om���AA��9?*�cd�$V4���GVA�.h�xo��is��ek�"ޯB�/�I����ѻU�cᐐ�ž:A9��[��UJ��G�==��U��^�������|9����T- ������?�i$j���%��P����I��^�k�j�ɗ�#AqqqZ�3�g�k�d+����|�������Ņ	?����"-��mh�842r��o�G��Mg�|�m=�;*��L�/ ��:&��$�����ap�]�mA�8h��H1f��8�K��+���R�Kb�K��K(�Kցp��m���������,�ڨ�s�	������њ��sh�s��m�����R�ı�K�R(�*ڃ\�����Ԙ=QI�"��ڃ(=��e�.?'�$ǯ��	$u��#G&E�A/	����eb��B#����&�� v�В7(޴�\+3GS��Ln�����nWaB?��S~��h�c1�"Z� ������F���0.��W�(�'=��.�J^BGbm]~���LJ�R�)����迈n����N����L��J$�]R�༛|Y��	g���(�UWccݲ���m���k��%����tB��/�W�HBe���2(��(��:�*�X�<�xs��$]���r�xc��R��S�Hl�*֒n�9�~a>�?�jX����[�#ʔ��h]$b��2�i`Q�ixL8ʴ�rzS��Ԇj��7Rᆹp%�g"rG��5�n�_`�/Z%��v
��`���{d�	%�f��t�!N��i���U=R��s��vn���DJU�uЊ3�eZf�3���)�g�	�ڑ�"嗻��#�z��ѹm�<�÷q�cd��ziv\L��U�|�����F����?i@�$�TW��p�C� ̇�CA�z��%���X7M�t.�;M��HK
\P(
F��0'}�j�U/U/*n��Z��ˌ�8��$"��|y"-K]J���h�+�eR]�W����l�6��L:�8{�mϘ���!Mt�E�6��yV��u48Cf���T�g]#	he�u��نD�"�5�␪rSh�,j�cCW1/NQN�;[櫎U����
�?Ɔ�F� A#���)�N��ósǰ��5i��̆���ُ,��r����7L{ �U�Uԕ�Fka�`�A��R���pM� ��(p�������n������|p)��C�э�D�{�CV���cv����b! . ���
m��LpD��1D�������[i�r})]M��,��V`ӯ(a�.rd�1zm��:M�p��HV�|g���B$CS�R��uE�UM���D�%/��Ƨ�K���~qIǽ8B�BB��8)	�I<yi꧕���|�.��o�y��4Ŝ���r Q
���N�SW!�{�CF���
�-w�ǹ��Nu���#�@�J_��;����2�_l?F�	�t~@���������{)����������U#w�&W!��v �E���"Y�L���b$yn�==��so��1��KY&%)��V�}UL�)4G��M������w�����y�����-\��$��d�ո�(�n:)~�#�+�wɽBc�<g��8�9�@�s��:;&O�hj' S�9.L6�{T����8��#�O@K�fʦ)���@}�Kܳ҉�b7L�Tj�{��Ĳ�w��N�&_?D�Zun�?U�1�dt����RpG��h��2w$�Iy-���紉��dÊ��}'�I]�W��u��(P�1eqO{Ң��h����H�]9�%�"wId�A�t�h�Z�uE0�	J
�^�^�B�䠣>r��IFAE}'F�=��G��%:��>����=	ul��'��)�*L��e��7�a�6�H��Ɠ�2|�n�����������Ԙ���$g��6��?L<�=�����̻���,��%�%lr��� �y�Ov����f.<����g�Bt�v!�r�/-:��aP�U�z*E��P����`���6��8�,Oj]�DY�Q��~Q�d�~�p��Cl+*aY+
���T��s! ��r�p��p��N��{��Ö�-��g�5��'+Mt$N�&{�P��T�'Hp<"}���Y�P�3t��Wq�̴�!��j��������A�:]Srz�+B�e�D�X�EZ�lR�C��7g�Q��Ӿ�u�\ߞO���X�0���B�y����\�6��&��o��?�<�	��B�0srk!(��	�***�:r^]]��,����������u��� ''���s����(**ʗ���f�g�/�ǍM�-��O����B�w�fH�\k�J�)�Q��)!n�~�B�ar�V�����Tt���\�R��J u�>�ѷ���и��m+��U�+\r��u��Bo�}��s�3��Mф���/�khF��_���ޜ�>~�r���� ��H�j�d|U��7���iF�t�9�X� ���5R����-�!m���3fWo���87^��5��P*��>C���!�����ES�bA�j8�����/bsE�$'����X.\����?H���A��ɐ���Y�q�����ieњ���B�hS�CyS ~��Bhamng�_W9��%{W�h��ѭV����###�i�q�]��>y�������?�?�@��Ǖ�����C-�ɓ'���U���paa�����������A��������}��aVV��Ԕ��_ZZ���xDD��������ׯ���uuu���/˙���1�CEof�{d������1{���H�����wJ�!��\����H���ߵ\�;��/� �Q�ƥ��*Y�$�P]�-�8|ږ�sl�`�7p\E�����n�	���}���(Wj�lnbh4k�iT���]�(���9r,2tp���-`���g)u�����o�k�ڻ�IR�ԝy;آ4�o�B	�OE��ʨ;��ZZO�<.�$Ec;��v�i�����x9z22��s`���7;PJ1�vTĂ���]�{��T}�E��D�3��E�\�3}
��2�4o?�τ�]���L]?�A�����!͔n`!�$e�� o���s�i˰F~���л��񔫯R����_v���� x�{�Z�~��>7�����V��- ��X@�*,@�7�г7�ǽ.k!{��� b���؀���rΏ��UZ�J�q�BԊ$/~py�-���P�ƅ�0�">�$��ⳄZ��DZC����䛨�<z\X��Q��8��J�������Ib�AGfi��$W����[(�{�����'-Q����?��[N�F��� @A=�{O{Bt7W�%��К�3�u-Ѯ�4Nc����6�/���ƪVQ�a��5W�X[� I&��2�}�/��ĕ�7���m4�oz�X�D�ZR�nx1a�Ȁ�.�ל�&Jd��H3s's3sS/SG��3�+b�H��_�)?|Ҏ `���/��1�ZG�~�b��@l���0��fY����^���}���<g⚛�.6��Tr�k��o��k��K�Ә�;s�S&��>���������ccc�011qqqA�!�JPP­ \rr�__v�A�!���tBBB�kد6ȁ���������5���]�E7�N���^��|�u��ܝ������e��d�K鉍M��i���u�F�˂�'VQ�bEW���Q��a�wr���Y���
�1�מ�E3����*QJ�菕H4���s��Ӄz=xY�̵	%Py��twS[t�1�_�$��42e��/*� ��kq?���6�
%��6��,Whp,_�U^m:n����iy�8]}img�A=��G�c
}ڈJ�[NJǻ�=�+T5x��0�*\*�+�7:�F��U�(��3	����G+Q�JώW�c=l0[VW��
P4x)U5�����[Y���	�[�h&�޴�_��53v�2q4v1�3s1��T;�}\�����\M����&��O~\;B������2���*���ߩxۑ��X u��s�̶����k��̌ ��n��rs��ջ�k3��`m�����>��Ǘ��3�ڪ�r�-ɡ25���Yc���'�]�����Y�o��nLp�ŷ�eMu��c��%'�����2�T��2�⦱�̗��]�1�@*�7�ޮ�<��r���_<�F)R��
=O
t��u����u��O�<:r���l��˚E7d����K�|��ѷZ�=x$::�m4'*((�������BV��=8�ܻc�t|��o�x*�ێ1N�D��b8�7m5 ��$�����R���'����<��^/�����?'��jo	���.�YN�*��j����n�n�$'����Ωr=w���7	pf7���SS	��kwk&p��{\귊��3y/N�x���E�������%�*�!p����}��:C�*K�~"!)Ir��k���Z^N$S<����>69��H;K��^5�TU�	�L���l-;ϻ��)��||��w����4�����0�Խ3�Х���$������Rq�1T���ܹ{W�h���{�������{y|8��I8�k���߼�?��.�;�)\�������*J�&#y//��.`�
�*�����a�����|���s��^��0�U�X�C���L�;+k�Y����w	'�J|?ua��=ӣ:P���7m��n?�E�qy�v����U�����8�zP1����T�@��=�7�~��._�~�O_�6��E��D묞�[��f�9���<�\��m�� �QJ�!$�ʁb� ĿO /��cEi��C�F�$'gh�(	hBպ flM�����l�̺��"4�SL?����
>D���"F��4"�y"ećNEx��1/�=F���T�vZ!�}(�f˸�1m�Tr��`u�8�@Y�aF�NN@�޶]���(5K��@YU����I
ZDf�Ny"��!"qBte)��*�e����0y��@��:�fk�AZ�v	}Em.�m���"TLᵶD�Lش�X�0��#P�
/✭ D`.k�	���g�x��(E��(�\���ب����<��}�m�Ta"\��T?�x����><��m{{��G�L0�6��{k�-�v�B������55u�D�Tk������v��l�"e�8Z��:F��!�\�U\�@f�ȶ"���Z�UqS�DZ��T�MK�uJ�*��B�D�t@)�4ܷ8�6���]��/�-f/��FS�H�4j7��=��@H��*R�e
�?W����s���7W�?'�@����s "�u�<D��!�@d��J;!�ub2I��kr������s�Es)�H!T�q� 5ډ�SDjo<ꟿC��i$d��xY�����4h��s��Eu��`"��vr3�ܢO!������,��h�]u���ؾ`��Lo���)�g�Xh[������'���F�1��D�L�E�*S��}ގ�e�'���o�`�7��+|�)�IC>\�࣓}�Ի��w]�D���x�)���Љ�s����iK�@��uG~���wI�f�d�'?�i�N{�	XhR|4�oς <�vSB�����;b�K�ӕ+(�Y���fN��ЕŔ�?�tM�z]l7�cD�4�Ϛ��6�L���ת�w�zl��ϯ�fXN�x: ådz�BȀ��2����{���[���&6m����Pw�k�Ã"8�+�n�j�(�ŝ_��6�3�+��^�j�x[���%q�Z3C����\����r���������/!{�6BxzzB^BN����a�ptt����w�����A3:�%�7ɵ	AgIb�^3���7S�,��Gz{�|;#wi�� ~����9h6d1K;˄f���"�ҋ�a�Wm��"�hh���R�*z̨/ۙ��C>�CM���c�D�O��ry���?��H�X�J�m�sD��C�y1�d�����5,:4���#!�ŃQ�l� -⮶�%F��{$�w�#��U�X����b�u�δ�i��xdV��J,c�	�S�C9�~<���J� �cN0A~��\Yi��p��ޗ4B�}
�M�����(]Bt��k?j|5��A�ڗ���Ie���ߚ�����jW��r���m�m�s���#���a��j'ǺJ�eʗ������A��pU�B�[�� ����|��(�W`���Q��r���C����ǽ��ͦ�`d��\/��7��l�7���j60_��F�V��_�@l�AJ�5������*����y�5v�zӲIfQ"M�q7�٘�Nq�S)j��_p������)��P?��Y�a��{��^���9�cLO>�zCm�xe��:�p�v��1���L�Z��F������E�!���;��y
Lg�S�O��6�����`p
�t}���漵N�rZ��+�Apo8��t��Gh�=�Ds���R�m�"�7�r����[0��rI˃ ���6T�� n���N��"�8|�_^R�pZ+��$�*c]ލ� ����l~�׭X��/]  ��Cv�[�������3	Bh;Y�;7���ZO�o�M~F�{55<~�Q�bͧ)6al�q�J]VvNv��tg�@�����C���ڥ�76��0�w+Ɋ����/>]{��|r���e�������d�}�ތ��P�L�n�h��b�ծ�3�Q�cev����_�XR�`��\ܻ%�N�ě����2��`���L*Qf��+X����c��,{Wzܹ>�,Ar�d���_�\�W������oK�V�#[�!�;�C��*<�+rEr��QW���EPFW�Q!Ó^��	(d��)'|���-���²0��r����=�t&$�}eyɤ��`�Lh�T�>vB8��웮�9�,����d�s���Z�7�ħ6~�	N����5 �*�Z�S1���f�+���t�9�h�eȇ���B���&h�ۏ�<�����X�Z��̂���FA;A�#)^K|f��aЃ��9 '�۰��.�G
7� �����-�$�b�����uhD!�c�9�BA��a��Z#�(�$1S٥aA/��wS��f0`����+� ���(s��,A��P�Pv�h�1G%nd�7�.ԭt�K����!�����ݻw���������C�555!2����5��-�y�Őc��%D��s�?�_!���5�rp��y�~
�w��� ®��>D��H�ZZZQ��=�.�4�������������v�H����''_ƿ��������B��k9�|L�h ԟ�>�D �l�೫P��}���BWJ�ͪ���E�����%m���-g�'��~.[p�\R��Ar��g��W�I=�'v�|
�gP��:25L"��1m��e��l���2��[��;�~,�Z���%&.�Y~��B��p�C}�>	�A�w��-S�q��~�B�w�ߗOF ��ز<�?<Yn��5�����\�i<��LX��s�T��eoNyd�L]��C<t��wac3^Y�$9(�-��6}���s���|�L��f
�_�t�⛃��7��f-����3Z{�1�f̀���,����sYA]'W�=����x!����>�"�iD�� �ty�P��A�BA&�V'��`*ᖷ���=ɹ��ܡ�BC9:��-L�Vn�?�v��]D��;9����]�x�o	�e�^5�Ν����M5
X�KH&������,_�@��UPc|��U�Tm0�+�0�?'���w�vU��\R::P�B��#�e���Bc� �hmj���7CB�n�V���{�xr��,�Ϸ��_x�6P���I��r�љ'
d-�\�T=�3(
��äl3MW@B����{�Va��uZB�a��:�bт��=�œ�G�����
�׮�`w�kz6�㓍��o�g%�V/K�C�#�M��:?�}N��E���v��R�}�ǒ��	x�mSz�i�UjK@��̈3����I�����0�M�ȏ>�DK)Մ��}���I,�|]��P�w?���U
[�^n��w?n�`z.Ú w�y7�j0&�?E�]6(��)���~5a."���d�5XR#�J��XR�cjZl���z6�Z��֪1S����Y�E�Օ0y�H�;���p�<�^5o�d�t�5�=P_��V����&�ȣ��̙m��r����#�PK@��FY
аrl�}^xL���XϦ
Qϳ�[ls޸d��wå_ڊ�K�
��Á��uL����t�Hα�v��Sj�%#	 ��n��W����+��?%�Ի�4����t��R����M�I"�:����Z����i`�e��\AC^2�Y�ٿL�/����i�˒P��B�!$��)�u�T��K�P�k��H	���
7����\lhh�WdBGK8�_��WQ1ΥT�K�E�3L|��7,��G�����x���d[V�:�>����C-F���ד��EYR8���J�%8%T���qOl�p1�I9�}Su,P���0�$���I�W�k��������/�(qG��c���}��?~;y"��"&Tnf�o����^���J�^�}�����ٞC�1��%�-7�
�����Q�9/8ğ��2��|������3�?C"��(k\���QI�H��:����|�\q�B3��}}���[bt��_iU#� ���6�9*�/,`�'��h>��õ1K�=3���r5�@6�����G`(�Ԡw���%�i� L�]����0��R���. 
�3	�Wd��{�Պ3x��F��-��2����yCw�I.��m�X��r'��1�W�]�/ ����QE��MTq���Ct1v�4����޿z�P�Fü߭�6�A�s4�s/ㅻ�p7�MqEcY�������/3��I��j������d�W�I�~hk7=�K_�����7���[���
�r�L�	����!�{��瓝C�`RE�1��$�u��wC"E���r�)�(�}0Fx�=�������p���ds�<��?Gk"&8�2����:ƿ`.m��ưI�Y�2P� Gc,|^��,�P�yP,$O��'J"$�ʥE���+`S¿>����� ,n�Z���fm|4��mȿ>�������>r�>"&|WN�P���"a�w�c
dVŹ�2_�_#����Y�&�	J3������x����.d�﷏h$A*i�~��ys�.����7�Q������A��\�5$�˷Ej�"XO��ϱ"K�q{���|^��J�1])(�,^4a]�0�Y6�����4�˝K���A���
Q��_ ����X9����T���0B��BDGwv��Q�~�x�V�n Uw�4KS:��X������l��_3 �f�C�V�_�VL�
��d÷�{��M3��fo��S����f����Ek�$�z�\�Ң��u��0�CQp�i&��q࿹5��"�Ӂ��zH
:�<c���������V~����:� ���/�jÞ�w����"����!����|!]؎v��M$ ��R�[
BE����Njp��R ;I�zk
m,n��Cx�n�m$����LoQ{��Ϩ(���6����Hz�3X�J 81B�z;�����o���}�����wt%��1W+ɮv�7Ӂ��(ՇpP@s֮��r�>��fq�wxz��^$�m�H&^1�	�Vs.<�@�`Xǫ\W��I2tE����� 'h|�t	��;�%1�TG>r���ip���h�@ Sے��Ι�9���.��Ā���Vi�z�
�;'1�^@V�]:� ��9 ٣A�޳r�W�����8#�N������y*;�pF����+|}�I���\تl9Z�`oJ_��(ȿ�I>�2��ĺ�2��\ �l������!n\,B)��xyHc"��H}����q�>�z&�d_$���9�g�&?{��N�'�9�z�m}�-�X�����ȋw�!�~#�2�D<�z�GDX>ˏ���>��:h����!���I%�z�.���%���\Ѱ�Ѹ��͑(60�/� �2��M�P��8{k33;s;�[Sa��`v�����ׯ���@.*�9��+<��vZ�<=:>�;��ѣgk���)޻��pd�	���9/ԖhQ�hr`x��>!%���T۵������2Y`U�x(��,��f�j�T��:�T9,���~jR����
&�r�_}�B�7r2b+r�Ȳ���#'���nwx�bݩ�=������D ���E�Km�%�Y6`�7�l&<�ؿ��6v�w�Z9F8�>��H�Fto��V�-bS= 7�~��H��`����[;X���'�c<�	�]��ο��	�L���MV5�����4;b	��.��%�K�B�}&��Xp�JF��Q�xX0ODD
�Ys@x":��l�Z��1E�3&�I�k����z/!���\dsz��㓾f��A����{�>'|x�4vG�j���	Ŭ��	��Ԧ1;1����	���i��A�* j��M�B0!�Q[���Bg=f�Tn)+u���Y[��(���K�(�ƕ�F(i]��S�t�i!��cw�`#���>T�*�?z⾦��KX�����$��֊2������)���ՐǶ�Sq���P�@T�Ik����\ll��u2[d�	�lĊRg~�1G$��S�U�J=ԃgE+�jH����
���7:1%�&��J��c:��6�i�JEA��3YdI҂j���>}h�����۩]������Cۢ�׻���@�Æv��+
z�I��SR� |�^]��:��F�S��s�o5YxU�Ĭ�����@�{4�#rh����[��*A+���G�C�K8��O�N�A�Ze@��B���J�~���"�S�lY��S#��W�	���W����O�o���d�*��>�����������׻5�g@|�կ�_��$���������{Y���,u��^a�ףgh�FI��fcccee�PFvvv<<<	��KG=�U>�f_f6�\l(m���P<B�a�mP�:@jt�I�{�SA�7/�O�z�?��t��/�I�K�{y����3}��%jǇ��b�qR�o8#���a�7U�����;99Z;�]*����f�^W}r���������n��IlD���|���B����ЁC���3�?Bq����2����N}O�A̪��S������MgG3����qh�\�|h~��&��ojA�9:�Ʊw��*C*���GQQ�k��3F�?Na;�#&&�[��,�n��z�Ϥ��Jׯ,ihat��ܞ,���Gj��9~Ao�3v_R"���_�q!���9���_���� Q������oc��2�a t���T=^3g{UV�D�ͧy��:�OXo����$&f��h!e[��p!�}W����JlZ�L�����q���%h{��'���*B�C�5%�(��"��ߪ��Y��d(�1���vn?������3�u����Ҭ�)�����-�Wc��������z�S�q[����oG P �)�V'�3��kD���o�bK�΃�� V��BT`	]��&���csjQ* '���S�H�	�y �eN�w3�"��J����c"���?Pr�<��Y�~վ���1��TQ��1Ŋ�J��	Z�z�<��@���X���O���$n��g�VՕf����B�?�`"��Mo{�ʟ�C��(��� ����r�8MR}r�4> �;%]�H�H{d���k���ĒR�-3^��w2�vF�zz�u6�8"O��cU"�,a�x�����_@�Z�/:I�#����rづ@o�5�53�O>k��O��Uc�!Uݎ�����i:B~3�HT�a��R�H�*>�u��k��Q�]�>���stO�Y�ة�,��/�9?�_�+d`-]�oc��9�5Z���m}d�+�,J�B;���A�_:Y��7�:R�$=M�ע4y�{Z]�q�)��� 2G��[��٨�z?(Ti���Gp��	�캔U�,3��=B���b�^������� >��sp7wq�65�����y�q[�~);�(�U\�	��ng�B@��!�����H�[$l��;<A����o�"_Ykk�ǽ��^>��b�_����舫�p��@�� �"w�%R<;��a��H-�˦~U�s�
�E�>]n]n��d����U�oR򚿄CZ�9�A���H�K��Y�������?R� Q�a�� mX^:DV "8�*�w��;���Il��G3:�����뎢�"8Zj58l�a�G�q
?��L��J޿:P>��H�+y��p���;ɳ�%�_���&�U�����
�$2O�R���	�k������l\�ֈ�L�ýx� �Q�w��n����� b� Yy�J�a��A��G��n��_�NjU���� `��r}���M�q����ɗ>5$:x�*K�ז���?b�>���j���Eh���#��&@�	LN���+G�Qrh4�%�@��2&�������_���ܺ��2���jJ)�w ��F�_�_�r��UE�;�gN�Y@������c��ݞ��B�7���%�oܣ�D�7���oJg�q����M�ʝ~�p2O�o{�+?$���[��2#��r������ܐ�\���4�-���,�6��A �כ��a��*~~ 5ǜ1 �Ma�CcaК��l-���?IF�٢V͍�V3���l����%F?�7��6.#x��@��o;m�Ѷ�,�jyyo\��oO�����,nF���%��n�8�+���UfhE"��X��R(�xɑ���Z*�'މڨwP>��P�XM�D�%�(��G]MTU���6�.���qj����3����i��D��Za'+I���X	騭�1�b&���$��04����)��QWlӅ�H�nŃ���YO�쟾��W~R���*͛r^z^�6�ۆ�֓n2�ɱ��5�e��)Qu��}?J|f���.�/H��v���Y*x���ȃzn��)���W���T5���������Y#��8²�U�FL����=�C�W���_O95�[gZ��w��&⡾�+Q�����%��ǟ?��%�����k��Z6n���y�2vj�U_ˮ- �0sM;(�@/*�F���I�q		��s�B?6�J�
:!�}D"V���I�k�I�����{�ĉB����Y����{��fF�|G��F�y�-��M�Rt��Y���*��_���M�����,sʻ��bb����>u�W '�5Ɛ��|�ޞ�J�}x���H�q���$��y������ω*��9�>n\/�#6R�����F���z���(}|-�s����z��fD��?&���q�9�~e 9們�����T_�K��ӻ��B�k��6CTn�F��ISz�B���#墀Y�%>΃Q��܂^����/�?^�Q. �¹���0e�x�������mn��t����R�4��Kd���_�>ѵ���8��DIPN��w�O�����ټ%��&����O`g�`�/q�vO�+�'��w3�V=6e����+��L���#�so�?u�9u��z�[$6���#��}�ucꟛ���o�A���A(Bg�	`�WD l��[�������h�1��
˾@I��뫛"�ѯfHk�	o�5�Tw>l%��a�-�fZ͢����c���w�^�A[��[�ˤ�Ǡ]7���4���-�Y��J�Q�M@�*�ᆟ�L"��"C̪-�=Q:	�����#�	���2�`��aS���F�Jm�`�Lc��:ڴ�Z�M�z�{U<U��"�]f�&��3���d_���X}��,@6����s@��#��+�$;�vxf8��+\	xaw�`�6%E���0Ϝ���;O�L�
�"�ؓ~<��U�� ׆�g�J~�o�dF@=xy����E*��k�ޟ�(�	M���-]��WaF��v=���������r���:�{�#Ǧ�.�CU�k	��F�`|�=:KS�1+|_gJ+����V��<��W��U��.T����p�0L�"~v>H��˓Ï ����0z���J��PS0���_�u}z��X��Q�l�~�:&�9��P�#�-IC���
�c���<����hN11��{SDif��iP��x�C�O��~��9�e	GoR��� ��i�\�Cu��I����|E���rx�̀쫈�k�p������]u�%�B˿q�dA���|�����K�^�R��;*�dRr#��$�@J\.ʾ�Ea}����R��/�j��zY[�]%����U�̗w/�����g��Vlf�Ϲ3bRЅ�)Sw �{�K0�K/b�]�zЦybX�1Ŝ]�'�g>�f6����G� �jR(
���׾Ľ��*ɟ��gG�F
+6���⩡���ૼ�CY�M�'8���}(�P?$�V\�[���B�Ң2�BNnbR:~��y�{� q�WC�e7A�:��,1�,��tQX�i�s�HZw"C�rL�X�sF�@�6�	�IƼ�Ọ�+�d�N$}����2&�XA[��[7�7�
�*���&Et��*�gd�-�e�q�W���Х���ӭwA����OA��ic�����-eܴ������[�֕}���B��o����(<{��#�mH=�4}c�5l��Z�3:ԍ�`�ޯ�j8%Pi<u /@��P��(�.@���B}(����ϫ_��\���+�_Y��;Ti�_��AB�!�}@�� �1%J*��@�5�d��Dkt��]�`���)�t)��	����y�w���x�Gk�hhxr�r��s�5�y��L����^I�8F��V�Zl��h�r��_� �m��^`>*o��"��w�pK���r��T1?�g���� C�u�ROQ�x%WUvpI�KN5}��ԟa"��o�#���d+�K+�u=C"�J�;�F����<z�w�u�s�F?`��=����j����N���Q��
[�巰�ڳ��F��6����������ă�����+D���\�j8j��� ��sB�Օ�ƇY�p��F��J{���	°|�٥f���e�[y��
Y��K���R����0=�����ku���m,X�|�C�Om�����c����Fm|w��I�a���6�+�&����"��MT�8X^����Y[[�Q���^�$.��a=�H�a{4�����[_����B�tB;��<|ry�&�9v�>ط������1=�e��S���Y$�(09ZNe��P^CŊ���$���tv8+�)@�}�"�#�@���twÌD4̚T;-/(�a3oD�}�T�7�_P:5�����<vG�:��Y���̣�\�cso�6}	XSSӹ��r�6 �� 7C���6bH�I��.c�t����(���%��l��������)�zȥe�yS.��sP_�<O��ěm`������'_�<Bg��ʜm�<�2.�WC�x�Hx�:1��N�C艅綹����O> ~�q�k��|���f$n�����-o�H�N��3Oܜ��^����Jԛs�-�Uc^��z����	#�T�j�69���+�)�~Щ��L�����s�&!��$o�R��k�.��m�*H�_"���;�>��G\��"����We��u�̣�_C���D��@Y�e�������;�����W~,n��z��fe?^�\�:tx�%�Q�v
�ۜ�ݛ6ٗr��b�G�3�<�˷��2�����#4'u6��D@��`�xT��0�~��O����Ұ���ʳԓ�@��
����5�v[�Ȏ��G-�k��d�B�P	Jp< ?�`�W.��	6U7iB�_�-��l����zѥy���U�k9onkǯ<S
ـ�2h��E�������l��P{���,�n��']�����3 =����MkEݟ������pձ�`�P�:�=����dC_"�}tn�B���fv��sk�4y�>��h'��g�b�Q�!���ᝉ��{�F�<X0��I���X,{��T���W�"8���0ix��1 9�c�J�����+tp�>��[(�'l!�~@4�?��k�B111��
QS����aeeeutt��䮡 :����0��M���?|����AfG�?�r�I˂	c�u���0눢�g��4���:�/y~f�Y���q�V�K>���#
��-}F��khm�_����ߊ}5�/[����6�)	����E���#��%4�_�0:�R6X<,� �^�y�z�m7*۰�&~�o�H��.ᑬ����r-���UWO\��QTT��͛���������ϟ?oll��!_zZK~�cO	�v���(?rzw��z>���V�t������^&���&��ƫr|��s(��%.�ׯ�X�s��Umk<(�o���kpݔ)#����W�b}�ʼ�1W�7cf���I!c�Ȳ%3R���h\���/��ѱ��>(�6^\�y]VlY�uޠ,���������]�l(��w�%nf&v����d�pU����tI	�����ه�MI�_��������s;�AY��8{�J3128 s}���J|j�X�A����bS.ٚD8)���4ې������8���,]��k- :� ��,��� ��%�'��@Ҹq�����7M��F�\.@H��A�Q��%	��Og����oBW/�f�WC��Qwkx�O�j�%f; P� j���0K�IM`�[�oN��0������?"�����(b^*oއN���ƿ1 �����\q�{
[3b<�B2�y#�yp��3�A��Уnm^�^{ć�.�OVXb`p�qV�����'>�er�;_�]���>�i��MW:-�f��55��>�=@e�W�J5b��%և�zef��q�W��])�3�C�7z�F(�����ə>H�Ț�-ӎ{/�������=t�	�	�@O���
i��~ig�����ʢ�\��ڏ�d�W>����Qַxz2׻u󂦝�#:=��3����&��֗�w�O�H���x8���h�K_zچ�3���4��\�zIF6J|��h�P¾ė)��q�����7D�)d�x�M7��O��?�m�������՝�Wm��b�۱C��/Ǯ�gI�6���K����FŲCWd�+���;�����Y^��]ϸ�^\t� y�7��v�����۲"{붜EFw��0y�����'��U�Z�Z�Y��p��P-y�Bnā�35(f�$Ի�Ve���6���*ͪ��~��N��M�O��.��������u,�$�o���dO�5�+c�ՙ[���D�ė4S��½�Æ��Y��yʠ3�މ���3t��K}�m��^h6��k���k��n�VIk�U:����Usۀ��t�a��ϐ�^A$�����%�n��[X��|l.
�ޛp�,`��UU��m������sg��h4��L�$Y�
\�!��4�I�g���$�=��@_tf@�j�?�� Fe���P����GB�dPY�X������]C��8~RP3~Yә���D�s=i3V�p��2��yJ�'����mf�ࣆa��|�>_r�Y�R�$���Ìi�^��eܦցtz����x%5{�gR�{>�	�����Yƾ��l�2�Kj�����VD������FIt ���$�����5�COo>�Aak�1i��n&�Z��Xь�+�Y���� �X�`@����yL�����`u3$��O���=��]I��?�F)�����m��NVwW���ֵC���H�����4�����p��;�Q�9�y��W��A�F�Q-�;��A���P.O���g����1N��~�}�Q�GF���9����V���}x%�iOY5ܔI5`4�_��}�x���jbEtWIR^9{O��M#fr3�_r\~���P՗)��14��q
�P�V�y)���{R���l��	�K|:Ғm���"� �X݋C���yg��,��S�AU����rg$��4֒���В[oq*�ͼ�5B��n�D %"�؃��ܓ2��d�c�PlM����cOBF�n6����߿�(���.�~=�	.Z���*D�Z���4���� �ӭ�J:D��ǯyv�0ާ9������`����/�GU2X)��͏
��<�.y��O~���Ts=M���	�!���|g*_[�(�����Sܒ,���1�B~��C���'�Lw�֗4BqNEkw(%
!)Wy-����@Y_
Ez��g���@+��e�+(�)")ĥI�L>��\�^`�y��˄\��,�4��O>�?ɫ��ϋB�{�}Q,֤�Qbv�Ŗ�>������q�md�5��^~�7\y:���c&ꥢ���`y&��S0�<1(�m L]���\�C�i��˰�8�*��)>�-�#lT��=�� ց�Y�a�2�V�-T;��6��������x��484�V>n�ǩ�)��:���"n�"�M.���B�K����`�掆�Zk�{FK=.�$����Qw�J��Ԧ��3\<_��K8�����'1��+�������1��S�S�D;4���H�S<`<.+���}#K���>��Yu﵇QlN�Oi���M)���v�e�K:�5��p�.�Ո;�5��߫��t?B����y�)J�Qb�<ʂA�`�\�!�H�8b{�X�`%�����S���É��qt6Fs�Բ�f��7*�u �w�)_;��VJhG�j�W����[5羵�OcK�"@sfѲu�^�-?��|�%Z }7��G�C�%�#8�YX8����Ξ��\);��Wo_9��~�.7����C�]�B��3�yڄ�'Q�c�Em�����	^�E�dE+�D����<����+�k�Q���VT�����:����E�G�4]��N|�7O�F>ݹ�25�9�u��������)���e�(C�N��͊%n��p1�7��+�"=��A�����@
z)���Ux���VM5!�:`��Ź�ʷ3��!/Ň�(7���Fr�����3���A/e��[�.:��H�u�~�I��mO���Hw	eΊM"�.J�Q'K���Bý�QR^���B������Z?2��pI޵�gT�1�������r߂�i7q��4ՠ�RŨY�Z�b�4�4�1���)nGi�zE$~~3���"���*�1�% ͆� XZ��<KV�}�n�l�S`��$��ur(��hs���G,�����eԧ���CIJK����]��$����4��������T��4��d����̸�����T��d��d��d���'9�>���O���}sӼs����oH
�j���J��,�ЗA�' DH?\��|!���h3�O 3�V:���S��iQ��
��E �*�\�7��_�T���� t�A o$ut�	V����J!��< �!@Q=����f�>��M�7o\�SS$xx�TZX^�lj4^�D&Y�G|J������Q�u�u#5�_h$Єkt��<�QO��2�1I �E�����S�S#^�l��(�Ú�sوA�_!i�`�=bl�߈��+�!G���1�k+�1hRk���hk�sO� ֘�W��َ1:>)9E�Ȍ��)%</<

�����4/�](�N���m�GkF�ܨ�826Q�V��T308��S����R\w���S"�!ipt��?6��?����߄�Lm%�@��_��!S�s�16��D,�0�ǄJ�aA�:���%dd��e��H&:F�h����h��-l�D�'�<�1IM���v��U�z"w�����Ղa�#��4��E�r�dj>�U��(j��(��X��c8���w�u�c^�C"�˲����4?�`w�_�
���m���2���Br��2�+�ap��)�T~��s���84�����|h�H��?�:=#�:�-�;2�WΣH�1�WM˕>豞v�Zh8m�z�(�3H�,�e=���Js�%��l�GX{��`%Z�p`a;���)/nm���1(x��e�����M�.�1�!D��і�� �������ł���(D%�4εꏜi���đ-p���"�/WEL�E`2��3_)�,��0^5��n	��s'�� �P�|�\�ש�޴�jb�O�1���1��1�0#���)�Q�Q����c3��>�wJ��2Цց \a�gv%���:���(I��#r8j�\����8{�9����ݠP��馮�K�$!H�M�����D/ o�����M���(V/�+�F�>��
y��8��_ �����C�y���?�[+�����N��d��K�u3ldX>f�c{���l��P�Q�mz��Bڃ��JUw�װPi��m{��J���v�hÇ�mKk��;�?��?�|D����f���W����y|�y��T]��4�	i� �hQ���Zc���L�Hj~�d�R*_��,3w:Ooż�u�B��v9N.)�o�]5 ��u�L���eIT������n��\� 
g�{.0�cIw��mS l%D?EjȨXh��cp��3M��4@@4��9>����>!�AH����<i�r��#���Q��j��
�R�H����uRO~����@�$�i9<���w���g濱�����_*���2�D�J��p�I��&���Q1l�����eM`-ӺE��ffIƪLvC�@���S�ǒ���׍��Ҹ�ƛJ��0�7#�Yİ}�Y���:�N��`D��
F���u�Q������{���gcwNY�=��A֯ԝ�l��g����rs�=��e9�Y~;���~��{8+9
�11z@|T�� �� 
8N�$F.4?k�c�O��o#L R*�Pf������)��|J-���j>�ㄶF_�@/`�b������
wooC}�ݷ�S"�O��>�lDk`��{�-A�?sZi��(x��`1#X ȅ�D��ݰϾ��j�@���c|�7� Ï���!j�`7��[�WY�������wն�)9��$O5��Z=�o����}'I61�b�3>�R�\�̄M���ն�\у1%�c�쫆UG:��p��+kË�C�3Y�v���3M#���4����뉏��}�{���t���u�؋��l{�o��d#|NG/>ou��A�D�%"":nA�vM͒�I`X�_X��ˈ��r�r��i��S����#0hO
	��:�(��^zi�8�k��0�­H�~��L� y8(6V��È�6�,>,�t�=/��f��R�SԱh�$���7�~�f1�>tus����K��0ѨeZ���M7�1�Ċ��Oy�����h��� h
9k�Hg��2�έi��X�{? ���A�"?VD�w&�{%^�`&:B_��/�a UN-�o�����j:������G8b�pv�'���u�
�w/��Y*��BM?������(
lf�f���N�����[g~?���{#f@F�s�/gZ�0'����8��E��9�L��j&����38u��)�'gI���9h�X_��D�d����O�b�`���?��O���E�D�}2�Fg�%wQ�d<'��gk��f�c�_"l��9�v���z58�_�-I�M5� ��
B����4��X>��c��ܟM�\�QV,o�6�h�p������R�Zt1��o�|��?	�5U�K~��8�į$�V"a����
*��@,	1�85 ��V��Bi�b��q��Px���LN��5��?����|��Ò�k��ZoF˄/7L_i�$�0����}��N>�S�f�CyS���}�b�: ���Go�m��s�%p� �4��j>,�X�(4U��=E	!�ձ��)TF��*x��_[q�tT �CK�XU��>�7�ݹi���		���SZ�A@ZiI����������|�s����=���}�Y��Z,��s�1�s�1�7	�@�7D,�V� +ԏ�R��/�^��t=?���Y��J���V�Z��S�;449���J�t��>7)�%t�sG�s�k
�W�9��Z�տ�m7����V�Չ�h)+2��ݝ2)��_5Hv��E����8��~)@e�IV}�Xr��he�D��fU�n�#���&�4m���3\2p!�N'��v��z��T@�ƇDq��<~)M�{^��Is���ö��yK����&Ëţ����bp���Z���A���|^���OCmY֙�n
`�h��s�BWT�e�&{�{J��cԡ�T��W4�kli��+(V|�l���a/��a�A��`���P#?ƺVu��Ρp:���6W��8ϴ@kj��M_-���î���f�����>�
�4�����?�M�$}Lx�Ѽb_v?��7H �ŕ���@�3�����w�;��TM8!žU_����f���bKע_���V/�|i�xZA�d[Zi���5�[��)ǆ�<HG0���SA�2��S7�U�#��y6.�O_B�h�#:��H�����A{��ü��k֯��Tԫ�Qv�����3Y�������'�qɏ4�b���s��x��������
D��6���=.��By
�S��P�?qd���Ke�/��f��#�5nFG)_��^�rI8[ ��L��^O��*�������L����]~�Nf$�<|�pF���9(�ުEH��6�Ba���D1��yL�D�&�!-��	a�2#��T��֦{'��O��@���W�,^м�/7D� �A�(|%�oxm��%b?܏���Y�������91���X����÷��	Rx�S���IN� �9�k�t���ի���?p|v���TO��#��
��)L����=,�y�.�<�t�3��ؒ�B�
=�����t���]cg�L�"�+�ĕG���}A���H����0�ȴpM���~�W��{a*Ľ�0ht��H��eJ%P��B�
��~~d�$��m��~L����滐�?�o��Cڝ�Ho�%�7h�2/�(�g�����z!�����Iƃ-�0�׃Hې�o8�Dp^꫘ꩦ���W����a; ��_=�>Dl��r=�Ჸ����1���O�R�d~_ Z$]͠їI>��d���r^����{b��G�f����}�Ki�ٜ,A^{�@4%:T�XE����-�������̑l�񛦺�2S��@J]]ݣ�j��!��?��U^ń�rq�ԃ��.L��a3/��+f
s�>yqܲ��1��͊:�,zw#��s��_���g�0�:Ml�c��,�is���^���O�D�� �?U5&���6�J�4�r�ذ�䇂�7����B�xH0��z�IUS7�2��xV�Z?���j$S�3��hk�IS���@����`�X��	��%b�ˈ�5@�H��Z(����,�<��d��a&����VZ�c����3�HĀ2�I��dF�',�Ph�~v�do�:S��[@K��z񺗃�l\zyBC���ٿm�����=���v��c3,<��	Oê�0����;�$�~b��Z����"�(�-�� �@������c�0�슪T,%6�Źs%%�6��ߐ����;�7᾿�����|ۋ~Q#�?�=4�/�C��'�  �����GσĨ%�>I~�Q��0= svɑ\���-�t�K$��<:��+�E_�3=O�����Lˌk'w����MXT'u��j��}����� �+��݅C	�d�Ŋ�Y��^�AQ~U԰ڪ��qw��<\+lY|Rc�r�v��d�U�R�Q�{~���TR�!%�� �C�|m^/�N�PJ��w<;Z�(ʷ�C_��K��_r��Y���{%�Hd�Uj��Xr���C(r4���*����vX���*��:Fha�QInM�"�R�l=\!��m�j�{���X����-�`�*
��:�O1��{�o�B��e��3�-f����F$jCFig���ojYni�_a����afW=P��k�i���D�<}I� �u��W��p䈐W�iF?3>$ė�������bǓ�\�o�-�-D�/ �~�O������BwY�>2=�=[MMMiii)))���BMM�ٳg����H4rl��K����s:9�p B�jM��`τz��	��ە@��0 �����}���$硺�\�dz^��s�����P�!�ގPcQ��Ca5M{ǴpP��]Y�S]��TP���/����	������� Z����4��12��)`�׃%ϟ��l
�-��4��cr�\�,��`F�XY���z����'c����*�1�� � �p�84��5�p8���[��t�0��/�B�O�1�:|e1��A�~P���ra�Q�c��A8�9�)N��`�Q�zA�X����*.8GJ���{t�����>���������D�M�g2~�H�\H�<x)i��qБm��%��V<�5|,�B|/� �d9�J�8H=��j:|x���tl��S�}���r+�`T��i�P����v�d3�&Bn��!D$�>Aك�.�O�����J��?�V��4cA�g��u�K��	�z޻���(??_4��r?h) G,�`�K,�J#Z$��*h�wͬX�:h�He7�\[U��5_��k�}�x��r�ȉ�|��u%q�x2���֚V�a�!?���A��8"
ۻ̦EP���8�Y��[�ae��O�DÇR��͉�Gg1����'{x�(Q� ��\���W�+���>����
���K͋/Cna��ZZrǔU(?s���5R(hD�;�f u '����-�M�8\�@���e�q����DJ�ib�3��JvT��x��	�/;��R)��E���j����%�?e������C�?�����Dz��E<ʕ���@<Jz���b��nRCaŔl��������q�Z���z���0�f
>�|�h۬�#/4,� �d����^7��K��'jqA��-�� d��0;��L\S#�&���}/��/�����V�.掆f�� rgI�z��hHJJjhh��?(k~���4���C(��/0h�����$L Tu v̍B%�&CK�Z�N������)�5(݆-؅3N<[[�M�P��I�mVBRz�v���WW�j�;gi�����_�}��m�E�~~=z��D2�iL��/My	��3���2ݜ������d��T�_/}%6z����7�F��K��!�W*<����? ��Ó�+�����'2�ۘL')�� d��z$��K�K~n�քd����VO��~=�_�m9��9j
ZE��'�K`�-�gD�M�Y�`>�
l�@����1zvs��0�&NVV��nll��d�6I�ϙx+ذ�cql���		���"p�] ��PjRR�n|Of�J�4[�L�85:>q%&�Ղ��$��;��2޻2���Pu3c_ֻ�h��鬕<'���؅y,11XI���VQ����2�y<=Юe���	���4���\�S�h ���"�c/܅���ł�R4 &�)���Z'ğ��O�����D#e�I&=����f�i�}T@k|=
�-.�'�	�P�iL�L%��oV��I0�z]u-ɋ�q�j�+*$`�o�aO�;LF3�wj��-W�5��6P�p��;M~Ţ��$��*�2ί�J��+eƱ~�H����TO���gUjEj���<HEm_�T��khhKl��G:�����]�c	Eq= &���_�����w���3��ֲ`%w�B�|�W��qv &�S�[q�6�Z�Z.���o@���b%�5b���6�7Pj���z5���=�&mY�)�չ5�,YSG
��K�~�RN��-���L�3��Ɓ�8�&fv������t��4ZL%�h̜(���z3٭��B�T w�/ٺ�a�b�^<��7�\_U#1����Fa�N���ֶ�<���e�0��&{��������_W>��16��J������8E�B;��z�݉�����;������/T�Ys%��t8$[�d�#�ȥ���E����q�2�8�p�ֹb'Y?��q�y�`� l{��4����aO{ �C �.O<��)u-bV��Y0���ؙ
-��,�P�摎�����h�D�"�%M!+�B�!���D�����eHg(������D�/CB��c��e��s��]Rb�:�?${���w�G�?�ϝ�-mm�nM��0"Ɲ���I���Y�P����[�.P_�9��!jQ�c3Z�t2L�(�O�<��h��Sw]�e��Xu>.\Q�m� @�S)
�����-ŭT���3�)��e~ٔ<ٖ<� �hd~Fl���1�Z�C_�������vFihl��MX�?+�2��;�5�R⾎��'vyu C=AD��j�Yl�wW_QE�GX#h�In!�G���a��t�o��Y��#Y�8�+�c	#S6z~����e1�����JH��F�<�vl|?\��/$
������Y׻=B���_�+O���m�����Ǡhc)�
��	B�&]��y���>Ln<* ��`�@��0�m����)��[����$]�"4�"�*%cU�J�;�n�R@G�����K�H4߲�K?"2�5��<�jV�G�9��Hlئ���L�|�F��m��6 %dL�
�z��i���Xq�I8-�;������Q�e��]:/��G�[����:�HFEq�8��)��^�����mL�X(���M�B�}�9(�z1X*,��!���f�&��^���FY�{A�l�@���/C��"�}5Y���=|�Px�-Mӿ����Pa�d�ԹcH�)�����s̜��9\A�3�wǖ�A�koj�J�0�v}j�&&��}@��E	�I��6E�Bߢ�#��	t�����'{�G�*
8*7���������6D��iH63��Ȁ��v��w�A_w�/¶ڵ���/�w�+��Q�!����\���7m���ϒ���������������C__���ۛ���C?�[/�����7466��/~K�_R��%R{�4�^�����������>��kFm�m��ٝ���F�B}`�~�O�%�,>����ˤ��c>
�.�4�>�X��F����q����T9�;̿��CU0T�T�+a�fR+͇uU���y�B��=4p440��v��������������@��9�wRa��6�s��K�u?<g���N<����P������W@9����w���M�U���&��ד�[���;ʤPWL�ȗ�xPӫGL�~��q�UA:�.;��A�O?Q����SR=j�r��nDkm��H#���a��nZ�F��2(�^sdaP'�GsUbf��N*�R ��d;�]��Rb��B]����<�򀂗Ć�G��T.^	~�*,]썠�b�۳��c4>��|�4M�R/��XŹy6K�3��A{n�2~�T}����ӯ��߳7���T=vX�VybA�8	�7j�-��x99N1?��� c� ����b/Ca�1ps�� -UaL���'��j���hXi�`u�^����1�~/��W�c̪�t�ev�n���/	d����t�)d�"�٦�������e���U�d�_���(.�0�n�]��H�[���#�앯���$��xk�y���x��.S�@�e�y��]S�n��Y;Rܧ��(�g�p|g�q��Q��E�&,W��V6AD���j!K��^���L�<�M�d�����;x�d��`ˤW�h��Qn:=#ZHW��0ⓞ=������r���oB�G�m;�I�=?g5ۑ�2!��'i�-;���MNP+��Yk(B5�.`\��i@u����">1B�H��e��7�*�"_%o׃x�[T�]W����q�9r�
�����	0y�<�U���~E]M������1��fA2@Y�/5�H���Im����W��L�D+���o���0��B_�g� D�o�0S��G*��(=5\p3W6+\��b�,cϑsh�p��/Sbrx���a�R+̲�4�ј��}|�0����c���?��p���U�䵺����$k"9��jr	��#_$�.E�Hߘ:Pn��~��?���Vw��xX��q��K^��1(0I�Y�1�GJ�5��3��T#�7%�}�@�W������;��dE`���Q���PVq�D�Q�Z�]a�^1����H�*P:�b|�?8���o!f��������s#��F�^6��Hl	Ee>��l��)�N<�-D�R��*��yf�meE�n������Dq��n��)ʗ�E��w��+.d������32���R��R�p��R/�vJW1��_q��.gs:�[��#���aJ������Y�'<��-���v�E�ض�@j��Gɧ�\�A	���:3v=0!�vKC>|�bJC��.�N9"*���r�����+�	)������	X�
sO堄�3F���ɹՓs�s��ҩj,%������`PF�UmKE�\�5*���a~F�<u�o!�$� �;���I=����Z��ǟ�ə$?s�,4�<f�>f�RAcIyN��u� ׷�_�0-�d�2� *�8=���ያ��j>���_4��'H�B��R×R=�f����L��&��W��mi5���!-�%}��桋���ҟ?�&|�8>�2ǵV�, ??
�&�J����R��R��1)\q�p��pK��mv��B�p_�H�
�N�Ǜ�ZMW�����'L�ٺx��#�缶3ݨ�ά��E��r�tݒ�H_|J�vSi�8�t�_O��9Z[��T��c�(�y��Pr;.ȅ4�O��5b�3m'�n)P<�>!�~�HW��B�Qf��f�a��=zd�&��B�����}\}"� �!�<�O$�E�6�Q���\�0�T
�R	8�6����y_��ʶ!!wA�`Z�Ȉ�>D�1g�j�c'�%�W��t�
�%���Ԗ�W�P��5���6�
B���fk5ܟu�%>�J���������L��72��o�v����^��t������q�@��g�t���\gA�aF
��]�7�D&I��Մ��iG���B�U^{�N j����'�=@�
)�i�1h]���z `�x���t�{j|��0�<��`a|$���%����ez�{�W.�?��$�&��j�[ ѷ��%���,��'З��Az��_ 5O��,�_��)��ԇ�rF�:CP�|)��
ƪ�a�״��4����*$���G�6�=���jI>2n�8�R�[�1���������B̖P�/`l�3��淋���J�����@�@p��]�:!�lU��?*�t����$�׹7�2���ސ���,<@�����N�����vb��yqo9C&`��)]��)6�����!�6o����,���u�ā�j~.mⓨ����GV�*�CC۪|�z�m42�:��x��D�ĺG:L����&�.V�O����FDv�m�z%e�E!��5����Y6�W< ��}��1 �K��7<~�e���4f�=��n����O�Yn��5?��tY̸y�cֿHztz���i�x�O������~'Zﹸ_��O�)id T+=[�g�@��+�W�Gh��RWɳD��p�Oqѣ����^Y4��R��J��kނ�aE�||��@X��t�;=�/l���e+��s����/��uGH���ȉ_�A��Q��Qy
$�������3��̝��ݞ�Gjt�pk�v�	H�S��K�Σ���>�&���sx��9��/A ��q4Lr��{�;G^���0S�ٿ�`y�j"�`ڡ��JAz��(���PS(g_y���D�G�7x�x>2��16����7C�昀i�pC�����y�|'/��u)��{>Ic<��3C�������� �i7��L��=WX}�?�V�� ����^����ͱ)^xd1��yx��&��jI.�*J��b��ryd0������oCO�\w�C"[�&�KU�͚�������2�h��C���H�����GR���eF`�0[���E:��Ӂ�p&�-Լ����a�0þ8�$�05�/[��3�A"��<5 >dC��#�X>%<�r���X�����`�J��q�a	}QS��7\�vp� _C³�KoBs�}������w��x��?@�MB�*mEڂ( ��W���]�����+��6�D��-�i��l����ohkH�H3�����f>ԣ8=uSX�҄�̈��^�&	���s��cdDU?hə�P#��8�<��fG����7�z�Ď=̰f�gO�<B.��u���P�������K����Y|2�a7�sנ���|L?8���.y���a7�-��������C
���5�9ݧ@�YF�w)!�|8d7(�IǛ��	�N�9��޵��K��N �9����9J9Ѩ�x�a�r���'&s�͉-��~���N��W�$�}(�p/��r��j��9�r���F+�]�kĆ��{ؑ�E��m��5�Sr�Kb��
�� >�깆����⋩!sޯ�:ZOI��ͪ�/sQ���ݪ�v�L�&5��
�I^<nL��H�|���)����sț�h�����mæ����׳�Y�S:�ϚO�_Lyl��].yM�T�
���;�V�?f�M&��V0	b卟�@�����
��-�!�1ƿlD�B��#r�N������4��?E��V�6֊ ��*7QNQi1<{$p!���&��Y��d��6�g 	2TB��iWR��Gq���Y���� ����ʷQ�v�B���d�ra7$ė���j䝥B�/�;�"�D	۟ ���y��E����dNq7<��{�-H� 
R0o����؛�OH�3^��[A�_Y��?�	B'M\1Б�I(q���H���vx2��yXg���x��A��8%��ⴣ�W�ޘ��o��'�9n��2�d�;m�l���-�k� �P�u�oH���0�eAU�Qc5�1���g�}^���� ��Ios$K4hh8�M(h�Cu(�EǇ��K]�~��#�_�����	��?x|l�����N	>y�!�B*���-<6��2j�}�2c=Ǚ�����?w�GEx&hd��*���=.v~~�|&������ۮF���������́��O�p��Dggg��V9����m%;���}�����]��@B��rrr:ng[~�vA�v��WU�f�2�(�|�Yj�4��^�C�$�r��~=v���8
�U[U&��c<�"�n;����W�B�L�ﵩ��Rt���,gST�[eٓ�!�a�}D�_�O9�mT�4���È�,J3=7'�i�Q G-�1(�w�5���)�Y������pG��Q��q:(��� RRRu�,��Ʃ��G��@�a�,+O8G�<
�;��I�:�+���t.e��=���o�'�����H�b����G���#D��5|��i�iZ֟�|��Z��2?�:;:��o����8\�rus�}��M�h<�'|;�C8~��)�$&����1(5�Noy��eor���\z�'��M1����/^\'B�y=���^��H4iy� ��CQ�c�D�R����G]�҃oDF×{	����hE9��᧘ Ayf���+3lv�Z)ű
�]p���-�s�c_0u\�\�SQ�m`o7�6;���bߐ;��3D�r',܈��b�;��|�PyyIx��B��Si]��������;77����&I!�������\z�N�77����ڥ���f �[3 ���'4BOWm6hZ��āS���H�O|jO�� �Yt�`����O}��Kn �}��3ȅ�`�Ԝ��$j�۷2����,�B�v��>��l�Y]K$������q��ۥp;�0��-O<g8	k�GVグ��^��a�I))�W�<!2I!NT�P���[o�������{&�o|ƅ$�=��:Hf�s��,�A�ª���V��P���iB�l���Ih�Y�H��3� JnM����0~NT�&�[�1ڼ��L� �^qמ�f�
�$��)�2���r'��� F��lK���=*�Ui�,�ߞ�4��>���m1PH�t�����}	�����K�7Q��;�S-��d�j�'����C�X��t+��ۤ��� z�,��	r�/���j�}�%��������@٨���'��CI|��[��]� )����0��^o��]�� �-��4�m�k�:Z7��K��f9���.&8�CXH�W�EL�
'{$V���O����雧����놇`|���
cu��`��bA��N)	6��>���l��5��u.Z�������R�_�k��!�
-=$I� �¼L�[�[%�M_�)3D�*�Y������&�}��h�*�fѫӜ����C�A�<i��^j6�|"�/��|c&Z&��z�-1[	5�f��⁐���������R��F���L�!tL�{� �����<e�݋����M
M����z��l����=�̨@]h~J7ն��'�}�|�I�_