F�4
iQ�^��f0�!�d]C;!��`���ΤS����@���4G:��L�e��6��� �4���{S4�H�Ƌ7�N�~�I=��w��j���hk�
��qY4��݀.��	�C��k��~�F+è������l#�p��������N���R	d����^�M���I/?kR���W��|�a�+�E��Fb��Zk!��L4�b���/�t�1i�^�� ~9
}t�����=��:�"�B���WL��&����v������)Bn+��V�oF)vP�m�6�"f3��$�̻�Go����^A�FbŚ�<��*�T�H�H���~�1������G��5�A�+6lI�fU���M��:����5yؤ������o��X���m����;��M��6��bޱ�倚�Ү�X?jxϷ�H�o�,
5��x��Φu���ĘMl_2n/�۱��Z��d7���m�¤w;e=X8غ�k�p�ܡ��r>�b��h�YԖ�_�L��k�͋~�8ce�V�_87��G�
,|< ��_�ίX�����R�k��tb��N�����r�W��L�8�����8�w�r�:o0�-�H�䖍vB�1�	��>m�i�=�Ec_�d�����l��$^Et����[A�XȂ�RM�EW־$�+5���b���R�Fy�z����[����,�{t��P�f/�Oʘ�������0��|_��ɯ��W�6�^�@'�v �u�U��a�g�Z+,1��t�5�i6�6�"�L�4	�N���YY�6��m2rد�2me�W���|��7���_�e߅�l�����m�^'�w5�K���_��o��(�Ə�}��#�y��6d��l�J�}{��q�H�ߊ��'��ZMc�GѨ�**?)b�����ѱ�g��S\�E�Tҡ�Я�`Q�	�8�Ц��n��_���ګx�̜�h�cq�+n����XN�h�$��Y�Ʊ�� +�"��O�(����q\7�@�
�y��B��V�\>j(���8�.Ө:�f ��,�.��og�i��] H�,��ٟ��9��:��U�|�S,�|*�����֜fQ�NW��/B5��h~���p}o,�r�Ģ���t"��Ne�B0S�]gb=�)G��!��OELU��it�e��[d���>{ʛf��I]%�(�����OO�蕳-�9������E�α(5���:ע����?���EO^ �9�\�;kD�mE��9d���֧83o��Ȣ� �o��s�K�Y�z����"����=�V�X4	���Rpc��JZ����c���ow��;W�آ*@|��S��r��چI��N@�0�ƥ 5�Z�̶���F�Y4�2�-*.�����,����� �1w�L���2ݘ�Y�!����T��0d��!��O,k��0�dU?rY3h���
hx�R�#���SM���{�ܕ-Y��= �"_|�E��K١�b(�/R�O�[�d�"GoKb�įSy�Г�h�k��:@��R���c^�ш���v��ޢi��rA%�����7VXt0���m#VZt��W�Y���'�(+�0���OC<��Ng�)��hk�\c(��I��RH˛���`�����x���*!�WbT.1 n|��_�ڢ�:W��c�j�Xt@��3?�x���Z����!��� ~�?�X�W����94�9��3�iߠ+xbJ�Ǆ���I$rͱ��h����slY�E���=^���?��]�g�(E����-t�y��<z����g�+ +�6���_?�yi�E�f?����,������~����Y����_��S������E?`��3���sq�E;s�jiL��bѭ[r�ji��բ�[s�ji|���^���',م6�yvar[ŝ������`oz��ݷ=wZ��n�>���m7T���W����7��>��Tŉ;=���E��}�}��������5<�3���-���Ai���ۏ���c�׼)��>W�q9�������l0�2��@��[����