C��O�h:��˛�ku��z�Q\�̀�w�LR��E���H()vq����F�Fm�Jj��LL��h�Y����nRd*RmO�_/ ��4��O-���KB�u�����6i+�����ʎA$���v��$qQ屡�|�
8V�����5;�����NueſN�87���8��uIBT/��.�WU(ܖRt���ĺ�w���.���WZq�ٺ��`�1��l_��*;�4��\I�<}P���'��������lqd�*�{��k��n0�5�gq��ǭd���u^�����s�5���ָ�q�'���&�ؓ9��:&��|SԬݺ�1�Y�L^9�oCaK�����,�ɧ�KR�f�g��]x˵�~U5$��� ��/e��Me�E_)��ݯ����/ިa�� �+�,���a������)��b)|�j+��~�l��MHDU�pR��:�eaG�ET6;��o{ԓxZ�O�h�"̠��R��E{��U��K�!R�L��7}fG-x;��{/��(5���f�٥,�b����=q��ݴq���ᆕ��fW,�����TÒe�#gC�\��+�-�?n�ɐ��*u����k�"��3�}0k���zf���6[ߤ�������D�3C
Z����2�S��ۡa�N��f��$e���d��_��&�8:{�z��~�����G�w���xw�&��H5���CܲܲYV�!���t�)9\)!pu-�n4tъ���f�S(�Zb��C� ��s
ڍd���&���7B9y9��{�˓��*�*��ٱa�����'`��q�{�o6�W���W�&ҘҘ4ÎӒ��| �E"5��V�iq����P���.�	��[�oI����~�4s%>�����@0�ܻ�0�x��t�
ˁR)6s�c�N�_��
����R\�kQ���5�x�bnfmJ�K{�'>�+��K�7�E����4�;��<bv�a�Ň�{c���6�`b�9"5��
?����w������Ϥ#b��^��}hcz�b"�	X���"l~��q���k�'>��_�W�<&�bQ��a~�*�eZ�;��^�p}~yR�+1r �đ�����)���}	�aw ���w"�豫{_�����y��M��T�(�%h(�U����lӇ*���O��z�Z���V�f:v�	�����<��3c�4�e��Zl�Εc��r�:�kx�B`�'i>��Eo��9�����8#b��]��k<p57Mf��������Ω��,��3��'侚)�1�/ �vĭ��a��)�WR,'�騎��A�AG)��r���d���v�c`��