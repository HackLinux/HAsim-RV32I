��s58��As� Tr�A�,%��Ƨ�P ��bP_��s �#~�s�s�,ͱ�As�s,,8"  T\~�1FF_<rP\%Tb�T5rs�,A�\s
] " sPrI�88s5
",NA�< \\,A%P?\rI _<N_�A_��PFNz��)s#�_�\,����,,1�1 ̑FFb%��,A�#�_,<�# ~���,A���rNr5 s˱N �I /���5,����P<���,��,�<#� "���A_<��  �ssssF�r  sI�<)F),Ɲ_ 55/T�8\�\N�A%�8 8]"5�"8�I""555A_?#�sP?NN \%,�_, _<I_�I�Fz<�~�\)�%P�<�<�)<#&F�F-�5A�\r�?�_\A<��#,r,�ٝrNNAI�5��A I,zN�,I ��˧_\N�� "s��N�,)�]������F�� ��99A_sٱ,I��I,,�N,��5A�s �"5r�\\]��" "�T\ %\/"P,z,<&AsTA,5 5, ,)?PN\A,P�,,#FN#~�,��<_�,N䙌� �?,-j�#F�9N!Ts���?#,\Nv9�-v,z��PA��ANr�z<��r_9)<��\r5s_���s
����PNA5�]����s_�����11_,�/��A_A#<N�\r�5<,�Ơ"s8"/�\,%8s�%8]// 
5T �55�� \\r, 
%%) ,? 
%%,#<)A,,#P??\_rA� _�<NN#z�_~<<�Nj~~��N��z,F�1z,�#&_�,�]�z,,<\99\F1-_zj1,_)�s~zv9z)s<�15NF�],���ˌ\s�r,#�~#A�� �r��%j����FF-?8�  �5AsA Arrr]b�
A��%��<,,5PI�s]T%�)]s ��\�/ / ,8 "55##< I#<Pr #AP,P� ��N_��,� s�_,N�<\P�z��z�ˌ�P  �sz1NP__�)�#��˵?N, �\)9_1N1)-1�N,\#�)v9,�P, \,sP\���"s����N��r]NN1F&�%����z��FFF�&) "]s�)��\%%�]�� \ #N��,r,)�r,�"   T\/s\rr�8A�

�" 
 
5,IP sAA<,<\#<_Ir#˗\sAs�P�\A#� Ar�̧̗���j< 
͌F���r��IN�_�,��,#)�_F_FF1--)NP,j�~_,
IA<5 �"]˗A
_�_�_N�����N�5��r�� #_�rN_5 / ��5�%�], 
!����
8�̌�N-1)P,,5!� "
�/%���s s�8/8  " TA 8
,\%A r %)ƌ# ,]�A,<Ar_�\���A#�s�I#\s\5I�ߗ�P����, <����P��ٗ��rAN����\#F�v91))P�zz<#!AA�r%,  s��PIr_\��#_��,sr)��ٱsT< ��
8���]
_,s���ˌ��)_z_--�#���AA5P%s�T��T�55�b] "T%% #%Ar#5 s�% ��~APsP�,,,<�s~��sIs��A~#�
P�z�s����sr���� ,N_����ss���#s�r� \�91#-)��?#,_b]�Ʊ�##%58��
�\ / �� Is_#r<P�\s��v,,s̝5
���IT
#j,_�A�~�A�NvjN�!�I�/,�8\s�����,ss]AN#s��rIT_/%## ]5_����s�<#�I P_��r,\PArrN�,�
5�AP�P��_,ss\s�ٱ_�#AAA�_� ,,��,˵_z_FF9)) \�)j&�\s�익��,#,
,)
�AI �)��%N�,A�s#&?_
�8s�N��\I�I��%%#,AA  ��ٝ��N!  j-̱
8%%,Is%%%����% � 5" s\r�A��
9_-)I,,�Ɨss,5,II~ss�Ň#s~__r<N_5�N s�˗���sr�NP���ٱ��P�r ,,�\�̗z��?sr/<NN_#P5<A�?A�P�s_�#�" ]_�%�\I/���_s,P�PN,N)_,TP&s �#-1�N<�5TI%5�~��NF��F, �=�P#
� \I\\�,5�5��,s~I5I\%,I8 8I5%s\P�)N=F)
#1& rs��r<<#A,����F#N_A_,A,N�,���#/�r��짌P��\#N�˗��  �5r�P\�Nz��z�?P\As_P5b,A��sAP,, % 555]�\�Fs�P\_&j�_z?�z1_~ /)-�?�_��
Tr%

88� F�zN��ّ�_\s8%�P\s��]�\8%%Ƨ<~)bb%"]!8\"88!  F1-)%]�\
  N%r���N�#�s��]#_�5!���AIPƱ���NA_�˗���Pz� �P�P��_NsP��zz_-&11,! T�
�%%N��N�,r  ?%
T~,#8�s��r88sP,ssA1v~_%P��\I�]"%%5)1jF�_���&~r�I "8I�I�s!�bT\%s�5)s_,\AAN//  )##I5_<,<sP_\,�_~_ ~�\�%%s�,)~���P�ˌ,]��z_��&��s��A\\�N��?,�z���F-j 
TI#9zv&N~, ,,A) <#)#�%r#��AA,�#\��-\N�z1��I �5\����Fj̝N�F&-&,A_\���~�%��5sPr5 5A5,N�P_,�5�#N
\ ,_,#,5%I\APA��s��rI�%
%

��A짠,�%\sA�s�z������,�r��?,)Fzz���FF1F  , 
"��F199<s�,,I,P,,##,N � �\_,,P�A,s s #�P\\1zNNrߧ%�� )-A�����)�)��F1N11FNr� ���I]�%5 <�A,"%,,PI8\��PN� 
 ,)_ PA5% rI, \��N\_�IP�P�IN#rI�%A�,#]��F�],�,䝵̌A_�\#����?,A_zN1NF�_~�N�

��˙_1F)19)��PI sr<j,,P�N�sr 