	����\�; o�/�&�����Þ�F�]�`��S���0�g>)����,��1C����=l%?e���*�)ǌ��<�vһ�	�T������ α�ulr	�W��|�z~Ѳ����J�R��Ė�^���dB�����e>!��m�:ң�/
��n�_"#u�rQw=�����Ps����{չ�e��蕭a,l
�Y���7�{���Q�/�`�9�7�=���W�˒J���#�؀��|�?&<mq%������~~�%�8���w_5j9�r�m�^?��0m���"����'P� ����xGd�A5�
#�c��*���@Ỳ��3���J�9�<O���Ui��ӳ�.|�.M�:�KNbŁذ�Fbw���Z���r�0�OE/j1��u�0�9Y�v���o����s���R��[�"��ӗ�吣W<y�-(�5��rZna�qj`3���ֱ0�F%�(�.��)C�ٕ�)���i�:�����X>������8jfu
���q��ͲS�Y�HGʥ���vm��}le��+�gB�$:sc��4l����l�jSIš����yr����\3fM{����f|�8-��I��%�q�e���*��ʍ�h��N������� u�"�k���j������+%�<�J;W��w\�V�M�Ϧ�{}LtJ�`�S��6_O����s�jc��W+�7�l����7�[��v�l�έ���R��9�y�ζ�$$�V+�l�vF�cDc�ޯ�dؼ��6�fq��v��;����5u
�����)�騿��2W�wK��]u�2���Fa�*r����l�_A�����z�i�k��[r�r����M�mm^�ZF!yr����Տa��\�9�&��҂������T��Wpy��iU]�u��\�p�� �`	�s�<�kf�,h^����kV,�>�G�w�Jj��,^~��E�L1�%!|�ꏅ���1������K:�$�p�ZQ���ֺ~�S������C�������?����p�է���g���0�y����R���իg���3���m�#�I��"��sN������s������>��^�hR�j��v�fE�?�����F=���j�Q,C�_����_v�g u�}2���V�)���ܼrd�sC��}�{���J_�O"93����R���/�@��F�/��k�%~M�:�C�Z�3�k�[��_J�)��
(��Om����#5�0��t\���8��<�Wb�����@	����i۩lP�I��ℵx%p&+mQ��g���T'�.�;&����-f�53��UE�����rT��=�CI�����'⧙I����u���#NV5����?)#:�{�����y#�l1[��~���̌)� ���i�tۂ�����q�����j�&_�c�	1K��""�K�_�b~P�`� U�X�<]�F�{}���v���+�?�ztx�X(�{ńz?����@�v�p���ƁS�ކQ
ȁ"l�<F��
*�@v{%U���y��1��!ٷQ�������K}��w�HhҕNW9��
G��8������P��.!ޘx�2q>Y���/���L���DO�k�_�M��>Ǉ���WW11�ϒ���D�8Z7�i�=K�_�N'����a4�o1��*��1�SSj3���1�o�װ68������Jk�����e�K��I�<���׶�JH�]����9��מ;����>`�8�A>̄��}=0t߱>pPP�IǺ1p}�R�7HH����U�$4)*-�¡,���)�W3_�ڬ�"A)7=ؘv0��y����������:f?~���v�>�d�t��'��Rr���-��k}9+����<�̓��xg����w�1M+�����*�u�Jc���-^�lh�ַ1}8z6���3�q�̈́�m0{F3�q����שP�}n}��x�]�&����_���˰U�!�|��w3��W������ft�������f[��ī����/�ɇ�F�Kڽ��t��u�c�f?d����n�����jjPPrYٺl�����o�I����e����a��<����r�{C���`\����j��|�Ku�\���7�ר]������t7���� ����b��w�J��;��^�������Tz��tq�<w�s|��F��mW��y/{q����t�Ԛ�Se��?�BY�"\jM� ��W�C��YO${���)D&��B,n��O,�.����Mv��Y����{F�95�6d��B�[��6�ZK6����{�L�q��۩=�/���r�� ���,�(N� ���'�	������v���T�YI#O9�ʇ2��^Dw������i�Qp��U�ƚ����Wc'�kG���CyǶ�u��ۢN�cG�n���W�g����O�N�e�]�%y���d�����έ����L��S��l�UG���8s��\6ZQ�	
��H�?/����G�Q��x�6U�_gTn".�֋�U���+���5WY�_������uFk��Cad����}4ק�XU�t#-n��[�����V����Ėd}�n&;-��g\��y�7w�s���x��8/���f�jnO@?�����<�m�BX��Y����`orv��֢�����M-���#�(n<�gT��h,(�-N�"������1�W��	ى�a=y�9���v��c�u����e��.Ϯ˼�ʯ�ۻ������-��I�Ӌ��l/Zw��QQL��q�l<��.�>�Dqo�ߵ�8Л]?V�B�ވ��;z��aݴ����ɪ�<���s}c�����r�뾑5����n}����櫑�Ka"��mk��X��Ά!�:c8��zHٚb���˲>���n�Թ=A:�A�	+{3��N��z3y��z����4�:7?눡0>�o��fo�6��zýҢ����!?)�bmXfukN����8B$�� �>%�{��>��n�6;�������4y���������K���v�k��4�l+�{�+�좟}'給֗�n'����~�Qgw��J7n�!�����y@Ӧ���psV�YV�F6�������-�#���p�}u�`dr~��A\���h�=����B���s=��a7[6��"V��n3� �@?�r�~�M�'pa��q���&��e����۳��lty�&t�'8�q1�d��{�y���a�=g
���Dަ�p9`�Ͼ�s�L��+7��
V���t���K�[��y��bѡ�$	]���nuK�X3V	z����b��������1���P��T�N|h��[�N��;zz���W����ь>/����	���b���p[���>�\OcT��\��+��V5eB�b<D���������̚1�@>B�R�PEg�/tON'����dQ��b�!%ޮz�Ԝ�$ޮ�Rd�+���*�x�bM-M;WN��?����t��I��'λ.q�����9�2�,��
�4z6ά�@�+��Й��
����]b�	HEk�f�������L6����I6SL\��!p��)��"&�zyԨ�苸��T��e	9׈gL�o˪l��/��e��B:��k�!�N5�u=[&�Ь(Z�h:�T՛g>Hq"b7r�`�f��w�|wJ��>����H5�b��.�3ݒ����.�����'t���}ڇ���}�C�u�|��w��m�H�v3��(�J�E����!ͧƼE�y�|WiS/jW�������!ǈ;����Ы�\K��軡,0��W�8���
t5��ex�@kX�Ё��9G6a�ɮ��-ʩg���m��v�B�T��%�������R��u�����kx�4n��YY`��������`+�hS�UF�Ί>�p�U��S��͟����D=u.���WS䈛�'�ȝ�c,i����D�M��\ʹ���6ؤ�'3���K�Z�t�h�U��"UV��f�mG�����c7���5���A�}6�+�y��C�c
��7�7��f�g�m�#��F��-JC��a*F���L^Ki��9Q�D`����B� )Q;���L̫B=C���<��L<a�u�ޖR������7�[�����B)$d��Ѣ��WSp�H�T}��ۑ��X�����^�:�o����4ɟM.��c��uA��T�wߤ�ƷT� ���ڜ�3��lZ��VS�!��q��U��r������㓵�;�æ���R?w���XW1s��S���� � j�r��G�����Ca����xJ-�г�R�@|3�����>��p�p�j@w��|߯�U�
���t!0�y���{�;}F���\�!d.�"��Y��gw�@ ��w�����~�@4�rQ1���ޕ��kJ1&�k艔�Em^mK�w����j�L��l�T�9�ˎ�D����p��|�f�����Lj�@���/��Z�'GD�/{w=Ti	)v:��|i�[0
�'���6�'}o��Dji�T*p�I?���h<��{ڳ�RM6i�ZbG�6�Q�Ά1.�Q�o��@R�A] 4`ߜה�b��y�>��77-��b�u���V[Z�HY���Ҩ��nje�{�gߐ����uѲ�p�j�Gqɋ+R�b&��ܼ<��J�G���� �K�>���o�d�8����5��^�j����WM������I�P�)��ǡR�"�$ת�,���FJ�db��Õ�{���K9��\�>�8���Z9�Ssy<�J4E��n���_�z�M���8��=�a��3lpWD��Y͗~m+���Z�����:t�U�=E[�v� ��!>~��.����m�9�3�RT�ac�ki\�r�?O�*��p�N�E����Ϊ�8Y�����SwƴM��e�Q{�|ƞM��Y��^��UN��Z�k��f��ܰ�J4�QnQe�e�/=�6�4ۢ�JoY�u�+�Z�=�k[Y��a%\�V2D�Q5D�:<K����$�ۉ����/�;?�6���:��jS�1jo��}���L�ܝU�-���2�,K+Tbt��Px3m��XC�X����2�dl=e��JT>g�C�L�~u���"��nA$������F21Ť�hcbIw{r�3|F4�M_{"�(F����������m��Ύ��3`��&sqc"(ac�B�=@>���J�p�� �{˰>��ˠ�g������e�	����+���t����EG��"�x�&7�����A��Bl99��u��<{D����6�UVߒ���7P��$O���l���?��#W�����G��?�c`�Ih
Ս9;����k~��Q�|��4�0���8;�4w=Y�NwȈ�!�����ҍ��-��͒xU�U�9��R�tPd�PdV�O?��K-��W���4���O�n��$d�:�[����{����wX�.7%�И�m�^������m8����@�,w܂aQYkz��!��n/FI�Ldk�����!;�:;�LFvMo����������8�GVïK5���V��3V���.�H�_/�YQq��0@��_b�G>l;KY��iZ�miz��"������Cf���*�t�ˢ 9�=���&��V����kK�����Gz�u�k&��*5�Z��H?�X�������ּ��ڔ�R��8�fW��,7�g��}�o���2-Z9�;��9�[)B���V�Ak/<h��#�"b�'F{gx�YΨ`K����N��}��ETT�e�[&ѐ���]��{U�|�����42=�;��z83R�!)�Ft"��f�� ��b��k���j�#)S��7�zT���f�g*�%|kXyY�'Tя���ӳ��Ġ�#�爨�{���o�{������$�.����Q4X����J��$��F���M�3�?�G�Z�Οo�<[|��/u��Du84�¿��'m���bcR�Q�cڂI� Jj�/�����>��-�S*a�
�QX�I�/�UyaXZV�P���h$���W����h���֎���G���,4�Ɠ��F�W�jdg���P��1��&��,|昣�n�}?�'�Y����M�ظ�����v�Y|f���fj|`������O�