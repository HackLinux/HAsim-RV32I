g�� w����T�{ڮ��3���mEp�F`"+�C��nl��F�/�������\#�Ҕo�h㼂|V�U(�����Se/�3CrL���wG?�aµ��>(�3&��r��ڼw#����ӱ��"�H�B$�=+&4��i���w��I��Q �"����q@��al/2xp�xz)Z�e�2$�i��td����e{���":��Ǡ2s� Zj������ݝ'�����D���
���j��'�W�>�C��L�%O�`A�?+$�����`��a�\}.���w�;�Go�=���gBL6@t�:m�������x�����ņ����X�z���AyN��ӄЙ���5����qd3��bh��M�.�o�.nq	�b�����|��Xo�Jr��k��]�=�`�/����H�ϕ�S�Kg0����A؝��2�v����n�n���
y�$���x%�~2�	� ������q�v"$�9֞�dH�n���i
³�znG�Y�v�az�7Gv� ,� ��}����g���G�����1�H��z����k�9��8���)��pxU
��������	�8,��46�jT�7m�_�g��&��(�x"@&�jl�)�`k�Z�@���fx
izh�%�q�4X+M��rr�3
�r��h���`��\J�2Q���K�,%���OPH�����0Ʃ��>`"g�,�e�S�]�+�+:���I�*}y�9{Th��L���_s�xBޚN�Ș~��/�$wv�Q���a=A� �a��4��aF���#���'��΋c� 6�vI��I{y״-�����ӣس~�Q@��?�ߪ�B;@t'wa��eO�G���T��z`aW,y�5�#Ӱ�2��߉�u��x�5�T�G � n�4e�q��괬������e���:[x(�%� rA��Mz;%8n���+��QX�ʳ�׷�q�Y@���W0��k�Ҩ�+�?7����������Y.u��!І��/��l�R�4������ ��Fߟ����������b�Ҹ�x��!�#~���[����/U��Ғ2���r�qp̄=�ZxX����,�a�D�?Q��$~�2B]p�)���L�6�X���wW��F��tPő�`W�P�zv`0	�n~�U=S���Q�l�E[)͐����N)��q���S�ð�C�s� '�V�i� VWx�K	�c���
�H�<�d��a|sy�<$uR�?X=;�*	������q ���jK�~O�z�r$K%�����
rt��#b�5Pm8�>���(��1>�����}�6�
X<�A����z.\t'�>�=>���MGf�}�������༣�Pg	@�E�,�9~���Dh�'q��ϸ�kYԡ�p���Ԗ}Dt�(�2.���jVMO��[ñ�70�yU��`K��55h�U��%��Y"���Q�	�G+���᝭���,B*i=���`xr�²tnG�󾅒R�`����T��oA%���L�I�B�c�"��6� �̿x�Q�T��)��zQ� ��9T���>�x��Q�r�)A�"-eux�ˀ낍�3yGj�A�{� ��Ҕ����$6�Q�YUy�	}��S�+�Q�뼤��o������Q��ok�25��;��)�9:}�x刞>T��Oߞb��+���D��'�/C�x2����1n):�z0���l�B��,`7[j��o��d��/�'g��G2@m�f1���|1�u��c��S�]�,�~�lh�O+qj�d�_��Q��C�%4�K��d��� ��>di&�5���^g�Ϡ�!w�S��R�6s�����4V�����h��J������l��4�1Z��(p�1��Y+pDd_2SyŠS��12�pq�����>��ސj�\��f�Q��O���"@�-��:/��:N�*`�W��s��Lc=tmU��q!�O�#��OP�=���_��rW����C�&v~ډR�DLn@�q�u��P*�hA��o�IKZ��o��J��\�#qn ����������G�ӚX*"����^7�Ԝ�����#Ri;���T���3�	��,G��N�Z'�3�aX[��6S��!��{\�𲼖�<�Q�����u�}�Д�,`�����8y:nfHO�J�"i�Y۲_f����L5�܇���Ph觠�p�X}�*��/*��9SG��ާH�ąIx%�V�>�~���+��k,��h��X��o���G >0�x&�ƓJS�x�PQu~t�?=B�V={E�
��f{���;����oV�!�i���|�� ���n�����^#�!�A��D+�Z�q������� �DT�Ǎ��Lc�Ƿ��?���T�t�����o�O e�gM�'��U5���a�0Jv��eX�n�i-lQ�~�m���H�m��0c�J���7j!�^A��u�r��22��i�.�H�� �@�A����-㛚|���8|dv�P�C0�k�o��kcK��8����3�����WG�Q��=V5d���>)�!��a��T$�Ӯu��κנT����&�x���D'3V?�r�'�aܵӭ�K2��M�!���]1hc��%KdU�΅q����<��N��pG�I�[>���c���V�|��q�J�R�Cʋ`w�P�ӭO)ˡ��9$gD� ��PL��CC�� h6����xu�K���"�"�fOE�5��I��iq��1�Gx�6%���������_e��n���J��~��l�SǶ�j��Z��sY��e�vڹ���4���ar�{��w��á:f�tR����C�	BAS�Y��]�^br����0f��zNyBٔ}|�wJc����=$ж�u�nH ��V�K��\�v?�m��X�p=�1�������j��+;�&�D�c���$á})5����	ͧ�Gj�D������vb1�'윸��D^a�&�P:�������C���|����Z�D��g��%�r@{"�S���(G�V�،���=���4��G�b.�^����؟ol#0��F��Z$�p"�>���dY��/�Ks>�($~��Mv����ƦSäʳ���}�	A��f�h����Q�?��.�|�$�<�����ݏ��1$2���w��6f�������`�8��r>m��`���* �j	�:�������v�Me�𪁣x-/��t���-T\��a�5�m���ww�=�_O�/�1vț�z�KCoXI�2�*��ʁ�,��UT�U�{ 9&f;����{wf�~Ur��ߋ�m��2f{������oz�`
!9���R%Θ,�y��l�|���X�H���S��Hg�
���lo���E�c.`�1��i�K����qG�HrU�g��Ir��G��h
>� �6�Ã����㬢+����Cb��2� �0u������e0�[�:t]�灊�J툃�N�+�V�w�'�J���}@�͓�_���`�>��Z��!a(��/��#�>�����B�kAvDW�,e�(۳X�j##U�_�loǞy�:##�=��b@ ˲8��2��+�SѢ;��}�����xM�b��)��u��f�"Io���B�����y��,	���V�*5\�'�&�i�X� ��8�#'�6W���5_e5�O2��*{��'J��:y0�  0�.�bz�T�����;�[�Mt@��T�[�ι��D�^!��9o���N	Q_|IX�DCБ�PY��s���n�����\(C*��~�B���QH��NW���I*!3\���I����2H-�N����J?�&ܪ�e�% 	F!��S"��n�>���oG�T��wr�8Q��..�/���BP)�x'��R���=�ݿɒq��wRں¦�X�X�cOs	�X=����ڷaN*�͵���%
4~��J���Plb��(�S�:�G�\��.�E�ټ�ԑ@P�Z�5��*n_��/٩�#�J8F�1�
�ƌ�h.�>S��ƬWTc����ٯy��Q׃E�=��o�ma�Du��=j�B��>���JLB¥
�����S/�5t8G�Bi�ۮ��O2���CVwgxj�s�������I�.��ݏ�K�\�m�M��_^P '�.8���՟��"5.��������e�d���o�7#�|h̀W��ϙG���9ΔiÏ�oOU	����eÙ|d����T�N���2�T@u���v���%�b6�r"c��A��,׃l�峭ޱ�c� ��p����l
{��+�����y���E�����U��n�*H�\G� i���n��j��pG.�m�-*��J�KW�bv��U����:��Ȗ3Mb�b���5���G��d����؈��¯�ۻuf���ȣ+"x����QTJ�d�Ao��@��)�p+,/fÇt��VL�p�B�(���i��U�4ì�^��ܴ�ֻ�,,�k�4�e�``n�s�aF7�7�#�b���p�7	�zx
��5�R ���$�L@ �k�o���|��Q8،c������[Q��7e?KJ9V�0mq�B�U��!�f/M�'��^,Qz��&��< �']�c���ה���]��}�5C괙e߹�v���{�IZÐ*{�I���Ju3��~X�%l�c����>��t2�����yE���H'�T�Ɣg�6���c��W���威�g�kV�V�<�&��������}?V`�����O�F� �2���eG�W��3.d�Tv3k�o<vP�ȅ�REdjR :�:'��8З+�y�`��^P�]c!.ՙ�!��z��@�C׺$�����,b���E"�3r�G�e����G�������v
�C�=��K�!T�s#7j96��w�$-��q�Z+�����0l)�I\2ȫ ��ʇ~���g��Y5� ��|u����|�a5��M�N�	E��A���s0��w֯�eǰt�G�G4�E�-C�ւ*�9�O�P"����� _�f�E�*dec~�[w����8#�Z������Y�P�<��4�ႢČ>��q���ƚxU�Yk�Z9A\�/]����yz���̌zuOfC�r.�����V�̘>x�*DA4
W�����W�ͪ+ �_��>�s�:�bl�ճ�8³V�l5�+�n���?��z�d@U�"����݌I����}T�nPbb��_3M`��<��fP���̭L�.6�/�S�*U���o�ѥ�Pɉe�m1&7����	xH%'�'�&�E��x�9F�t�ԷŅ1�c�5:��bΰ]���:]͕�ʒ"��b�b�M����K-ZR���м!�p���/@b2��({���N� ��QA�d�j�[���@�|g"v�~d�e�E��Y�_����AX�cpp�����P��=�+.:����/�w k�ϱ��@���g���/a2�K	p�1�鰫��-�_Ϙ�h�bJ��nH��|ɭ�x0y���������?���q?���*�Յ�����B��������A!�,E��+=�kRɄ}����
s���"\P�`*�H�)C9h��������󁂵��ﺅ<w|7~ɿ��L��9)	A��7(����w.~�r�%8�cG��g�ޅ����/��;��ߠ̒|	�Ǎ�5���k_�9��Ng�*/_�����4�
izy��uHv��A�h/�t�L%�9�=��a阄y����|\��� w602�K���6��g'x�t��y�2DD�`�Q��c<�H�~�i"�A���m�~$t��
(�\O��*�!t��������tȾH*gw������6�H�������ʱvX��F��Ȩd!������(-1��M��$�x
�>,��>Lb90���8��g���!Cn��f���^Yٽ�	zG	�|�E�R[n�A�T��Z�Z�b�wڴ���c��f@�g@7�K�k���\��2��ϊ���a������o��gg7�2�u�9�r}-���s޳���}Ώ��܎��P�oR�`� ��T��ѵ����'�U�|ऩ�1��G�8��R��Z3�ףa�eۦԉ��!�(�b�����NLn�ty��H�׭����:�q�Iw"��P!�+�)l��ٺ�����U�`Ec�,�p�Ǜ�G|�{�D��n}�kf@
�L��*�.n��f���W�#�U���UK�u��Up�c����d����B�'�eZ��t̲@B�v�{���늈���Lw�M�f6�DJGed�����;WV�K��YCX쳳3B�3��Z���0���7���D��H�=�<�m^Y�s*x�0lo�����Ї�)�-aK:�Oݼ�z��ţFD��aJⱚl��K�����a�I�{>����������~�H�م$�aC�FBcT;7b�����d�6275��Q�700e��0��/޷��k�j�ZDh�
�/n�4�݁(�}�~sLu�rT��'ؽ���N��z)g+'ċH���n|}��a�L֜e���%�1�(� a�֐nn�d��u�@AD@G���X����JNg�n��]3�~=�X�*UZa���Qx`�OYv���AAGK�z\g�na��m��'O<�٠�u�LJ��:��P�[�_�\d��?ݸ��<Wb��/�]��0ʊ�)�Nƃ.Zd50AB�@G�gO3ZG�O���V��	6.m�l1Q�����=uI���rM����y2���VO���|V����=�O�֣�65����E7!����|������;Z�"+߀�`�p��IB ����cL�{������������E��I2ҁ��)_L0���J3����JW%�K����L��C�T\�f�|}�I��f�����{WJ��w�zJ	�'CF��&l���v�Z!�sNX�T�D5WU��<��wu���FԿf�N>��#�2�2}�Z����t0`Ҍ�66���T=Kd�J�RP��4����x9y��5�f�-��Ԩ����.B��OC,6}={��0]gIcN���
�x2�����,:t�vu{�D�!/��&
�qN�G֡�f)�$X/p��o���ݝk̺�9��X�|Je���HӬ܂t/ﾖĖ�*rX��u�HL��>�$R����РEJ�ǀq��/���cPP�hv����ϰn�,��.}������]@���}v��e?�>R)<SX��2�3K��M_�[!6���G:1��vN�f���a���f�l��]�|I�w$CK	F��u�r��l��B�4�,�s�FU#^s<Œ4�X��k��Z#�����,¼�&�`͉�X�p�#ſtW٫#�
ȉ�v����j`.e���s��T�s�I�7m0e�'��u�XF�ek�>� �r(	w0~�
�ذ�'�N2�ڳ	�#T�R�M�p�a�`�/���u����`..D��1����L�����-ӫH��H���SPaG��RI�J��X$������S��5ɚ�hC)�h������G�rƲ��gC�Nu��,հ@}�FS���x���tΞ�ː9Z�ƔC�%���b�e�Ƃ.�I����hH����̇�sE}γw�4��G�Elc����[a�/�����hM�T��<���IGf�����X�{@M���������)�Ѫ]��ftnB=Q�\hiH�/�*Y�1�f�)B�����IJ�m��y%BI+H�I��{�O�v����s�u�L6� ��+��U/�<7�"~<���-��g�]�smE<�*`3��K��)��Y�a�yv)��O�"��҉llS��l38�8��8��l��
�C�N��f��(l�����L�*�g��i��]Rø5;t�hC�5�\���͎���L�읥�����-b ��a��J�?e��I����Z���_D3��U�|�̟a	��:���3`��t7���a��m)��:��ƬQ�����!���s7��� O�(@�G������=D�]���fd��q2��:.�;I�!�g�,c��F+,g�Nb�@�[(�z�����&�K.�@]��<���t��U��=wL�'Y�1)�-�`�J��,�;���*�gq�E5w6TL/O��|��(��(%��_�y�`���J��� _H�|�@`ގ�f�������g������&��"�a��!�L$@�dm�t�m;x\�L�Lte,^��Ǎ��<�IAݒK/%x��Ȩ̰U��1aK�V�!�����u�SItU���I���dK�s��,��Y��*V�x�A�[���[�2��|���P��w�6��g��3��K�j�B>��y�`f�t(��H"������Xܷaɣ3�r�)�o�I2cw�G��PM��7�w�j8x5w�X�쩕7��H������WJi�H�m'A�b�U�<QOoK#T�ڏ���
/B�p2쁹���Hr�`\����"���3�m�
��������I�1��1h���y5gl�[��`~�+j�h�f)������2��f���i�r&�7���h0�V<� ���g�k�]w����.D���j��[�,�u��=�V:���D�j=~_olŌ~�G�f��I���L��(��I"���M_�7I���f�0�م�O���_gd ;_�݀ω�F����i?�������0�^yH5C�T�<���*���{E����u���'h�A����(����t��k��K�o�I2�(̋����p7`�gB�����d��3��#q�ei/� ]�`d���$]�c*s�'nN�cW��B�s�
4�f�V?��4M�,��	v�[�D�g��WIӴ�Y��+��e��P�H(����oH�0n��F���JaA`Z���Oc��WI�q�"p�"�N$���I�x��+5U�a�Qm��p�a��J�Ѵz6'�� :C���6��h�K"��Q��Nnv�Ͷ���w����8�CN��N��b(�Z�37O���d�q��F�
G���`#���FΞ֢t�D�a
�Mgo���ԥ���e��e�,t���L��ʨ]�����d�M��5b��p�(�l��g5Dzk\�z�~Uۂ��*�:r�Y]r�E��[l5�2x���Q;��9Z���O�^rٜ��<� �r�TB����[��d��|��q��q���\���60�v��n
���p�>˞���ح�7�-�m�8dљ��ߑ$s1Q��"���37%V��1��$�׸����Jp�F6���MԢё��M��q0�'vޠd���Mt��@���]��u_u��x�f8�6NŇ-�ü8��} �.�ܒ#"ؒc�t[�5���Li+�x;���Dv<k��&����f@�#�5��iI�UM5��4��+���^ඔ^�l_����^V����FW`)8�"L�b�������"�m���Ӷ��6��u쮟=���>F ��������(-�Ӟ��	�\-�J���!D�=��\Xނ_X��]X�F�"�����P�Yc�<�KUlSoY��T�C��N:"ة�@<�rh����:���Yդ���\躒������8�X��� �g;��E?�P~�����"�� ��Z��y���+3A`;��g����vo�����ȇ����O~����ݞ��C��y�B�y�BJ�y`����R7Z�9�*���2�y`�7�ՌC��eގ
��q�XS�}�Ş#��<�=�%!�$!��j�L&��lm��Ĕ�t�B.�{��^���}D�X��ݸ@��J��b��Uf)�@R���=QG'v�c������5� �|�'[uB��sM������)�>�'/Q��^��gJ:9��;z�dTQ&"x�)~�WZ�UZ�:�osO�l9=�D9=ݤ9�7A��R����lO>�WT�9�	��j ���s�p�s�	�Nm���z�_T��_�멒t�m3�*J�bT_c�(
y��KWm�Y:f2����YѺ���ϟO˥��W����P,�74i|�l፤�h�hDt�*��iQ�ɤ�s�u��A�[�%?sM0��\c1�����Cl��3���J+��F+w�F���]A�8uC�KPx߁>d=���&�*��:�(q�w!��Pa�o�7��%p�9@������k{:�e�Sr�]���'��/'��o&����~>�ͱd���!�*`�	mw� zC��j>jܯއ��e��]!}z��R���}� ]��`no��f6�PĽԃ��j,�;l�p��(z���-Ƶ����҅����F�����b��|3om:��� �@���󿷙�Q�5�4x�h��0��~���ˇ��qlK�v��yѢ��G�������E�sx4:|%��9rc�t�1�Va�����~:lD\�����3L��C&kb����7@�֠�ǠŚ���Si�{���&j�ˍ�#z���=����9�#ֵ��Gݑ�������
�f��������&Ne�OJ�S��F_*��s�6�����hYć���t��nXã� ���o��j,�ޝ2����B�]������{�S��R�.�8~��U[U�R[U���d.3�4��l^.g����l9^�|�<��g)���u�I�4�,�5_��5_��]���6���6��<}Mk����5���5QBk�ʑ�ePkե�'���'9�rk��\�~��&>t��j�@�~jr.l�4�'[���5�+����������f�*������w�fZ�(WO�8��8`�%�>Z2�W�V�V�0 K9{R��CR�@���- *�=Ԍ�Y�6�`@����Y4L�Y4�鹉�������!�ѥ���l�֡�Ap��$���YB^����V�n�r�M��f�<��Es4�zW4��&œD�	j�Y����E��%����e3�ph3�tf|Ԛ'�W�����.�Mq|t�!jH��Nŉ�K�i�K�q�S,��&�?!�?ѻ�e���+w��l��]���,�;��AOfL��]�d_���@"��n �9GZ�C�Yf�>�{Ri�h��
�zpB���
c��� D\\rC�b~C���aL�k'�q�>���壤��{E���@����	���Y��AEb5ф�� �#��K�����v�$��������_�l����y�]ퟁjx��;��ds��;oX%��̩����c��]����J�����,lb�d�WjF�餕:�bA1�$d;����Jm!�-���2��m��t�ηZ�O�p�vh"j$�&V�e���Jc�������\bQ�L�(�t�unL]Šb`��i����'3�����߶��CZvc*��*
~!
>"
>��i��K^4�)
)C"
)�)
)� 
)�a:]۾:��:�ܛ�����ល��d:�&�f"��f��5m�˂����(������i��z�f�N�J#�������	��A�d.������!�{��B[�!$d*���z��
jl)F��)q'l˯��GӴ�H�<����<�q+r�E��'h̯bh����	�0�7��:D��h�=ŏ䚦��K���<m�<j-�}����4��-�}����]B!jx�n�L�����{a1��3�"ؤ��#��Fj��Ǣ�1Q��nvk�}H����f�����CjEy�'��߲P>mD9�/m�<���D����M���_�u2�ܔ����{�ɾ��KzX���B i�n�+荗��^��Ck{gߺ}��ܚ���a ��|B&SY4�s}ԥ���`%t#��ؽ���;�k$)����Am�$m�m�x���#�!��[b{%|�뛹L���`&~��
�!��j(s�x�S$jD )����Ud�Sn��������������������"-	f}͊$�$:��[�t�U��ݠ�� �I��>����H����WZ��3��\�Ւ�"�w9���U�n3�^���*�ʋs��H�>+i��ʕ�L�z�e�4��^�J�Ό�^��3�x�u	��L���Z�����2�⮹���H��Z����M��� [>n�t��4i�s�A\�"F(n��,�-�d�u�����,b. ���r�|b �B�=q����s��c�U����L6G�d6�u3+>�h�i�T��>�5���H��H�cf6�bp6�bT6yd;	�`5	�����������x-o�[��)҄��䈏�|��u�����kOEs8�&�ʼZ�v�;/�N�7�Ċ��k1����lf/!��/���aZ��*���y��ay��3���r���*�L�x̊�� Ҧ-i�`�So���-`�*�{��l���|����/����o1llJ��,}U�#h�E־%~+,���������Ʀ���Ɓ�������6e k�|���c�|��9������Ex��)��E��Y � ����"�����Nb���z����N���w&]���c3�J�$�tT�&�͗�sݨ�ʞ�ܸr;�a�˙l��ھ��l��e���ڹ�+�������iV[wk���$��tΘt�̻�V\�G%p`��ykۮA=�P������uÍu��u�M���:��t�-��V�l ֆ����A/(U�^���	���T_���y�_蜍3�F	����;xu%,���ÑkP\����a�z�2}���6���6���6�Y1(5�ԏ�,l�Q�T���*�(��V!��j!z�-�->g��k'0"gK���uσ�K���Hy�8���Uu�@:���y�<}�X��?���Rt܂��9<�}WZԄ�F*0B.>��u��;��lg}/����r���;�̶D�tq�4<p�7p�%p-��e]�eE֥=ya(�f;������}�{��["�[ES}[ƹ3���S.i?�!�@+���4�r7� �l>��荥W]��]�N��4� CS��-&��NI�+���s1��j�n1�^�O蚗H��WY��TY��%	�e�HuJS���IrK�P����˼�#/ݽH�&g&	�Uj},�B��{�ʻ:B�s?�k.��
�x�˿+G�E�]�)m�|b��G�ꑆ3���
�_�⟣gh:�8�E_�T-�����k]��X�RAi:���5�!��,����F��f ���B�Q�e֛}Y���'�5{	)(m[K���Cn:S0����i	` kb�ԙt�D;n��1rD��/���|��6sCa�ԙꨇ�3�h���'��E��E��u�M��z[0�'AE�sg�؜j�,m�(�����a��h뒶����������a����B�%�㗦�����)��癡6�����+��q�o�K���:�e�i�8F���E7l�=�����~"��K�-�q~�k�vlg&�㑧��N���k�7X��85���6e�W���t�(��vd���1ui+��k�����ÜKz�g�l����"� rB��;�F�C��!�����&��dֹ�X�C�#����jl��g���r��	���������t�y�_c%+���F�Ҩ6��!�q�3�w���q��Ϯ��ފ��6���g#�p0ޢ`���d�k*BE�󏍋����c�������m�o*kj�`�x3�x�h��T���������ǡ��/kbv��;�����zƦ��/l�9�531���j�V=��v����Cn�$i�fT+7/ȶ���ڠ@��efA�����Vz�-i,�g��(�־�60�x��g+I颂EV�e��U/�~�Р���1�/|��D��F��
s�aMo-y�V cg*���&i+i`�����;5�^��ir�V*�:B���?C3;F��?�	��5��$��A����Wug����W� ���G�zF��xFl�x�&�n������ %2
q��A���x�X4/������T}��xR�h��{Th�,\*:�s@�RV���Ѥ5Z.]LM���b@g����|�.�$"U�c
Z��$�M�h��E+t�|>pz=�ӄA5"�I!�ɉ�(���{�ԁ.����%#�S�}�ƅ|^���N��1�k�^����2F �!�2��O_4�E�EY���v�����#)��7���L凙��y
��įMp�����ֿ�'�?)F��'���'������M�]�9�dX��� ��eu������^��_ �e��� U�u�%�Ķ���-8�% q-�Q�"�;�̔�e-�>|�S߲�$L�� �����ÿ���N᭒���3s7��k�Kx-���#k��tV����g�����fkG�uK�Y�������$�����]d;n$�⤊���2���j��j�Z��M��=�NX�4.�IhL��h�z�`i� ,�m;�S��6����%������Ԭ���3�������G#cYi5���r;�`<��6Y�^��O��>���X�rB;��E;?���&Пw�X��n;Τ��J�n��An+5����n4a�i�}��^rl�@�ވ�Yh�Qa5�'*���G�kn5xv������by��й�d����;�d�f�!�����k����7K�YB���b/���&���c��ii�ai����T�E�p�`��/���[��=�������9�y��]�b-��Z�Ą�FſI幄�#����4O��F\.���3o�Ҩ�5A��K�5[G�H�۔����z����ȫ������iȤ��c:v��Y�Ϙ�t�-�M4XV�5XVw@���a=��,�d���x���X��bB�e㹞��U4�qu@���>uǦ
\���)��X��1��#`/��_��B�Aݰ^D,7�G�Y��^��!�S�AXn�9�����!!����>ɕ|-W'e-�~�~�5Z�7Z������"�7Z������F\�h�q���c��/�ٖ�,W>ݕ"p���/~wW\/�u�h�eH�ש/���G'j������k��ꈌ5�<���>:�sR(J=����L�5�3dP��]S��\�d��p�=�4	���S�)L�}L���ek�s�V�g�[]V'�!�I�O�㏕�Ƅ)O�:�R��U5���>��FW���_��%)MM�]�Dw��nʆ2��/9>�]�q�.��2��_	a>�S��B:�e�s��_�=O'r������(J<M����P�~�����<��m-��⇔(���}�g��/Fo���چ���U�7�Ky�h��(���-Iڿ�̆4�T����)�^�Wk����Z�4yܖJ�2��:�e�U�i����,�5A��zԗP	�%�U$
:�}�%{BB�����y�>98a�_., 'U.�wzv!�=��mޠg��%j�sY���G���������^l��o�Y�3�j����wc�$���а��Xܴ�}�g���1��է�8�52.Ӏ2��Z�Q�4ϻ��o��=mE0k�er�3.O�z#�~���ǧ���3H�OY|�-�S&�J�9���(�F���D��&U>���Q�~�R��*b�G��ʚ��}jx��(���g��F����PYoCMP�V	��e�+�'|u�}L��+��{��vc����qD�a:�N��J��o�N��Q-�{W�C�����Y<�{�jv����<���}r2"1��PjE�&3�<Ž�C���ONN���R�Bf�-���A���/�O �AOG1��*�3�2Ռ�2�:�`�*�$[��?oa�ף-��;ie�!?z��_ꝙ����v�fh�9.��0��u�*:P� �-Hd��&61{��tg���6j)�e��f{�)-�@�&���hd�-��ӌ�7m(H�`P�]���2�����q�;10��K���t�!U��,i��a�#�Et�-��=P�%CH�Ǒ���W�L����?�!yѡBB�1l�O�h�{Ew���N��$<�L`}���� {Ԝ8�=eq{���H�	<Tk�������my�u�I�|%��fE"���qW�̬�ߒ��,�EH0����.e�]:B!0eц@8�-V�i���x�3�Ke��5�w�7$��)�f�M ���?(��H�d�?}�*9 HQ��
������)2��|﷮���|���5j}C�G�H�{�#L ӛKE�7$���lSa�k�u������8�d�9��I��|�sHk�'�����Gb�Ga��,�B:�fm�d��qQO��S����z���C���l���R���{�&-a�.��97k�W�]��}~r��8�趔��J�����С�yW閪�}����O6�V{E%��&�:dևTԪ:d��뙴�H�w��Q�;}�q��M��3�m��H.^���*�<P��M.�"1�z���<��~��rV�~a�ׇ�~�-��Q�	j�z|��͎P���f��er�fa�9�
:���ş��u���g�@���[��£NtfQ^nD8��/�P��UQX��EY��-�M@��>�}��`�����N���Ƹ�7i|DL�����i���U<�:׏gQB��gH�Ѧ�@�Z�~7����!ގ���*�;�h}�7��-�Ϋ����!|lyD�n����h�_e�^G�f��y,�"R�z�#>`z�����`(�w�M�X�b�T�ڴx�x��A�Kg���
�h$ �� ~�ۛ�eGEw'zJ(Xa���vvJ���Q���s�i�`�zWo\Dp�:�K�Vc����!W�#�7�6#W���ۅ��,d$��%�f�X�T���4+�t�����1���vV���vM���)��	��ZY���������[ZRtӱV�H|"����5�-zS�Im��x��!�QO�|%M��{�7���NjMۆ�rvDVL�[�I-���a�B8���f'��H��iC��obu�fu,2���$�h^5#��ӳ�<��6�����P%KD�g�����J���!P��z��2����P����ӌ�WXhB�]�'fG�e|�x�+��Jc<��|��}�%�M#�`
\�$�&3��F��!z�;Ŧ���~҈(�z7s䬏�'��K��i�8H�+z��{����bp��V���ȳ��Ć��܈8���f�-�az.��ү�I��N��ПM� ���`t��l�;��0}%�(���35�9ݺx�rav?��<��v���Aש��^+� ф���eȺ�������9�Jc�gP�����������|��yW�(���>�������,��ǃ.�u�.J�e�6!���H��i�Y�]�5�x&l�'��I\�t�/X�"t$���Nx������JjL�5�D��Qh ��)N�}"(��w��|���i�,O�/)��[[Wh5�t����:f+�r�?(������ѡ�c�H�+4�B���R&�m����处o-�h�6�C�H$/ϗ����Tr����l���`Ĵi+�s�`�%�o�2�P{�Z�#��D�&�ʽ��H�|%�U$6����s̡���&��N�I�@1�x��(�I�5�u}V��0R�~~��_i�*��(��_��+���3C�K��|�sx�`����է��p+����ǅZD>��m�nB	M>��S"U:P:]�:��R5�? �Z�_^YX�l��Ed����5���γ�L���N�� .����F&���AHGFA@GF�ҕ�I�d�6���4������B׹�����چ�c�K�F��pͼ�v�6h���W�`$���2� �X7��n8r�st��T�f%�!�Vx��!^��r������~W��m`P$���N�.�%�ʝ�.ݔf@�w"sOD|���n�	��g��{�ݒl�L�gG�t��ۙ��w������V�n`�$��g"1U`m��~�r���lG�~��J���^N|��8�uN&���l����c�j���x=wtj��g�ķ�m��ﶘ.�a}���0~7����=X��6��lPѪS/{,ߔ�k:D5��w���`t�0�B�@��|�-:%�R$�!���v?�|����o����Zk���:�9NꗲJ�m��`�N�<i�W��m�R$�5�ar�r��z�H3��0�1�j�P��l�S#��oj�.Y��{3��+���Ok\�x������3(��5m�E@�'��J�d����?hBm����s)�D{,��6�Aq����H�Y�2��.�Dyل(�v�´/ҙ=$�P#�@`�(���츽���� ��d�x�,{,��Dٵ��l��M��T^H�'�szC�mp-rQ�ݬ������+���&x���������LMi��$��(���({�y�t� ��.٨��0&��ָh�������NZ��B2M�E$�����3���޳�3�Ǟ�  Ҷ�cT026�1�GDK@��C8��{z�+�������;��N)�ϚѶ���C�t�Ї��h�QW���GB@�4O�zO����G��7/\�.L�N�pj��O�'{CO
ֵŧ�dt����B�1�N#����Ѱ�]8�<�T�H f�ۂX.�#�s��OKHG�!���R�B�7� _c��P��.��²����F��^ex�G�2�H�Ґ�H6g����O��X�d��۩���xh�dQ����1����MEC �`��W�\�/ϱ0h��N��}J�Щ�~?=D�l�NP�L���l�ܝ>J���+��c���.[U�kJy��79�F����i($7������b�l{�IK�+�/���$����7"�%���7hC͚��͐o��U=`Nq�⢡|a~�����حi��J)Hd9����ay�T]�%��AB��*Ff��W��%�Ȏ�8ӛ�DF�9X� ��f��B%Q��U8��+���
�F��7v Ң,]�����זGy�?�N��G���ܷ0��k�h�ʍ��j�p����:���޹�·���h�U�+�V+�w���q�`z�㞋/�j;�I{�Pi�G`�S�SP��U(P$��"Z��b�2��ax\���񨷰�yxI�7��0I�9A�����ikk�)KK�K1�&��g��N�Q�V�0�*~�W,�?78�P�����7��_��Z�N�����|�n���`�b�8�y��]�x�j��߸ )}I9�[5���w����B�}i�ȡ5��iiv{����V�!ZII�0D���}mpHAA'��3�oqvi@~yð/�d�b�L��[��b2�V�ɂ�/smH�a��GO@����ž�TRղ�6��/�)*U�c*�6��e��栿�o�K��qs#|�V�y�1L��n�&��@Jj�7#�w�T�������Y���?T`�*,�7��x�0�o�+���r{ߨ	�+ыC!��ش��X~���?��⃑����IM\7��]D�1�NOL��詈�yK�Zf{�z�(0�hu�`�����oohAx���`�B������н�o��`5��42UC�wpw!�	n�;/��yߖ�s�(G^�	p	����C:`8��ӢF�h���ح2�IX�U_���J}��U��;�`��D1�`�����H�V��hE}$zk��ʯ8G�a�u1����x�5㱁�W鱊����}G�?�3Ty�T�,q�<�������6�k`���Q���GmO�ʎ��@�����I3���H�j�=:�Q!������E��Y8�,D��1�:jt��#������t�$jL���.j<f�s�q�9B��MOԏ�i��J|F�ۿ$�(Ӗ�7�^��zi<�?f!�c��!rn���֔?8��h1ё:~���f,�5��+`l��MyW�Z@���@ih��i�,6OG1�R����eO�9��KrA׭|��YK�	4�M��yzT�,��D��K�G���1�@h�)G���'SP�sPGyL��7��۾2V'��uKs**YM{	�3�(ӐF_�O�Mv`C�f�e�tɨz���G<��J���X�2])P�8+Bk�>FSw��X0I� �?�W�,���yDJ��G����&�|�D�(��t1� �BQGCw# �lvC������6�j72P x�(@(�U������~�O�6��:����&�g�R�ca[٩�
@�LN��Qh�V4>�"5��wR�e2��	�y5���<\�S����ݴC����;�q�
0���ۣu#�ab`�)r��e^�И����Ž'��s�($=���������[��1�r`�x�m�g�"��)vm�_t��V��:Y�.�_we�s��`H�R�(�&*�#��GefM?��P"F�똍���鄄	�l_�`��ޓ��VE���PW�Sw��~DfmY�T'Z8^�R��)Oc��H���9��
3���ψծ���	w����\W�i���Ѝus�N��0ӏ��'T��کn�V�{'�G�f�w�R+ .|Θv�O��vxpQ�3B�b��l�&t[�ǧ����)QХD�s�|/��s`�D3]dmc����@����·��Z�����I�C��)���!����9.2�L ��?Eu#��N�@x��n�AM�:��ų�ۗ.������gXO���x2�����9t(6K�>(��{�c_"4��� ��'gp~�����EP�|���ջ3��L�<�>��	ÞG@�7s�w�.#��G�M��R��N���4q�Y�����RB�ݬ���[p׺{FC�j�K[kJI��u�_��=��ߴ�"�X�#ռb�z��1�TaZ�Z�����(�%�n��`��MjYKT��-,hKڮ
���N�-T���LE�_<�5��֎���P8����o�}i'���*�J��X�:?���U�XV�o�}�L��aш�}Y��$7y�%OHk�k��f�#�-F��;�#��;V�.s����FK|!ܔ'H�BSYО�D �cE���<��JB�B�	�K��q�����>�[��e�A!<=6 -��,ӯTt
�s�_ya]�kI���:���}�4J�kݵG.�09�����bџ�$�9�������}�h��J(�)2��b���+N�h~(gڜ4����&:��]���:jtӷ�~�N�N}�sǅ,�g���SL1G8���嶫�K��l����w�V�ڠ�q.�CK��T����������B�� ��$���}�|�3�+����8$�j�Bpf,є`��*��sިw��yC��f�������)
P|`���ʆ�2�Ȃ��!Z�C�@!}]�w� ��Jx�c*'��l�dU�T���?NK�|�G׎�"	C�`���qNs�8����z1�_v�yƂNk�9����F%�����Ĩ與�qB˽6��M����'9�H�TM�T��=&?/���U�$@��DB|�$������gž� ���w2ԣt#u\�.�dP�_`Cj�;6��}����UCm��l	5�\f��e"ӓqy�{�O5��8.���C���6H�8���.\h��ǧ�3���U2Ӓ�I��N\ּ)n�����(����x.򠷵/�n
\>�%}K�����#k�NI�G3�u���(Q/po-ܑ.$���~������!!��:�X��zSW�9;�	iJ݌J�+���r���(&��)$]/�Y1,yb�P�l�Nr�w2�n�C�霟>eְ�1��P���K��<��4g���dC���{I��u ���]� �����V�[#>(I�څ@����a!_q�F9GhMzE]\?��I���]^IjCnu���k�6+��ML���T}9Էk.p�<����I�����m� ��{6X�g�3�
c���Ҷ�%��z(��Vv�����6[E�Yv�6���F�9��~LE	�s%���#2�A�Af�c�*O�d	0(�=:���W��9!����(T&�)����+�}+������KU�2I|�����Y"L��q=B���;y+�ם{��rV*�?깡˟�N��w����"5<Ђ����]�ۧ�?.L�;�s�n ]\��0,<�s�GJ�Pj����۸>O�M�P��<a�
�V�rr��%�ϡ�����,[Iщ��m\��L�ZUF�)9D���6��k���ߢ�R`=vH�������aD
:��$if����Ep��^��•�ޔ�Ӽ��έ�������%T���:�}7�*dCiP���I@U�Ci#�������� (��r�3x}q���j���y����J��	W�p\����xl���B=}\���FJZ�.[���;-��Fh����x�]/P���fn�������,�h$�Z6,��~_�Q佾_s<��]e�R_�D���q�1=����5�B0��S���m&{;�J�d����5t��@Dۇ��tr�-��`ӮK�y�d�D���x�V�m���ܬ���B�r�|����MAx���|� ��g�����*#s���s�	㳐j��E^�����0�����/����ĭ�����K��UK��X/�9���w��T6�17�SY�o�4��g�z����ַ�lPڤɊ�-��@n���π�Ɵ�f<��ē+�^��βT��[p<"��D8�		�~��s��w�Ĭd�A��$v$}n�g�R�(G�S�����?o%D�d�¬���!us@��3�}���4�#���wɣ�o��b�(���4�|�g3o��`�>�<��U@B���\:��*Ic�s��L�BE�%�;eŅ�������|�\�^\���5��3�����p�<&q��c�h$B�|HT�s�j����"�6�\a�ӻ������B�%A�s~�\�Ń��`�w ��9Fǎ�~�!n~VS�ѿ̶��ߣM�zF���"4K��Z���DTp���]�[d�*�R��g��I��D�s�D�>/�Q^ �U �_;��ө�������M~z�k�zт��(��`~{������t��jȱ������|�XW��a_#�@D��6��at��Sj��%��.�i֗�u���
i�G��tA��u�9xZ�yE+�OQn���9��3��݋�z��G�8c�2��+8+�+./p�8k�5RR���1�w���k�~eI�-l��]g{u�3���;���N?>U �ZtV�h-�
�Ĝ����VF��GP����?��z����4�B<�Bhx'tO���/zօ/67x��ڑ��I��@����:��P�ԭ-*/+Jg��-���Շ�xW�)�fCKD�t��({CֽT¿o�o@�+x��F|Ƒ�ϻ��ByQ��th:�gz�y]��C��$��&���)r��tI�xцj��s����\��1�V�~y*,���Ҽ�zv��8lӏ��`դ����iMT���z��r}!1x	���0KS������R���]��tT��(�������oIM���R���OK��=�۰e��e}8��"��E��_��$�q�1'<55-<'�+������#4��+���Ȭ[d�*�\Mjd��ȅ>����[��"��m�̯�b���S��)��P�p�g]i�¬�Wꎴ�G����U�g��F(2�I�*sw|�𑣕@��i��42�PP��n �e8t}ST����	�!;�n*�r��T=������&a.)+� �^b�����y���.�\IUJ���- \�f+fT�����Uo.4�s���r/z����,}IM�:��l�d��g���U�a8��Y�um4���ο]|���v|�yxV��s󇮾����f�>��t�/��U�Ft���uB~M�Y���^��(QW`n)���D;ȩ15d	�P�@���WX�yhl���g?�-�+p�>G|ƥ�¯������mc�?r�]�6Y��l�'6y�W�y��	��H�׀��{a�-��m�sr�ԉJ�Jh�-�:��h�OJ�o6�ب�{�j�ׇ.o�L@W�V�Nj_�G@U��ƲuN�G?y�l�����x%�����"w��œB��-{y���N�Do��1]�BgV�C����g��J�!��2��V]l��ɖ=2���|�ϑ�R�}�@�G�����0�r�t�hϥ�����S�ɢ��h/+l1:R�q���X/֍�
�Q�[~k�wDi�>���cs� ��OB����Mމ�u�ï.1���4="v�jֽ+j�_gp5�ֈR{�����f�����^%����܀k
7�����=�^$��5��hW"F`�!q	7}�ֺ*�p��U��Zc(��,�ЈT}�K"�h	S|��<�Ӑl���e�qF���f������S|��|�[�l�g~휔��k�f�J�}�j7��ÖMoM�f��eTe+����X"�7������l{�l@���l#`$ֈT}�	�`���
��jս+j7HG�U׺*M84�z�ѻ-�
9��{��5��
�^����2����Y����ݢ��Ў����4��>�+zmһ-������'jE�>����=��R���l�<���цو�����u�85���ӻ-ܜ8�����[l˚h��R{��s�I�m�`y�m���l�7����#m|#gP$����ީ��w�ax+�
L-����N��kZ~%aK"���Wد��q�g~�&�H��0@$�����N�jm�ax��߮c���`y2���h�q�g~'�V���x�2���\@��&�I��15L}0�N`��Ez�S|vO#l�C$=��������6����.�B�ax��L�����N`z���7�'4��B�\l�M$��T@��׳�պ*�=��z{��c����a�i�=�)��Ѽ,K.S`�;���=%��P��"�S|6l���3��Ѽ,k`��}2�)ֽ+J*^G��-�:$����!�*;��+�	\|���[*�7��
�B�*��f�<��($�6 be;+�5��ki�ّ޷:}�M���e;џ��s�����f��R-X�5��nh��nQF�虶�7� ���
[�,�V�5�5�8�&d}ihѲP�D�6
b���Y�&�����A0�֭*�F��qz�-J�q��k�t���A������qR%��8���!�.�wsdB壵�����c�>�j��]�.�;��
O&LPĦ��q�m�JE��l� ����8�#�����W���y�*�̀"���WX�5jm����0�����ut�B�b8�����ݟ�Ê�ĵ1�=�����`�=��q4S:��1G5����H�tvd�SW��kf�8�|��O�w�&�Fw�G0��k�X8E��u��%ERB��0"����N��+�%E��ٚ#jpaҝWC��a�(a�o�R�c����-�a,+������5ʸ�B����	�`��5C��U���6½r�v��N��h`��.�j�c�{��Lt����4�}ur��zЬ����Oۚ���(��&?�XCDtWm���7�	�<����V��1���!���T�����3�
T �_�A9m$�vxUo�p���FIH[��Ɠ��4,�`���AT	 D)�3�RԂV����_�wUp�Q�7O�\H ��|�6���j�T��lS~��c@�}�����7(dC�+���������h���1o���RAd�E"/,v�I�BG��7h���F+)�"�S��њ�@7�v���DEo2	B� ؋�Νu�d$�G�y�'�a��ph�`��XN�Jۡ�Ơ�/���ɩ�]Λk\����#Z3lV2%�)�w��8�����*F��з��!��湠�(^O�g2��X��LV1Ա�>!�������I.���N���P���CC@D_��U�A��ި���sSe+T���s �6וz��z^~"Rŋw����[��qt�S�p�xb���q�����؞����I �ܛ�i��,�M}_���FPp��P0���8.��-ܯ�2��@kґ�� �E��֚�����Ig
�����������B��2!�^��
0��xC|lO��x�l;3}�y3����I��N����	�!@ě	!_�����ŉ�}O�z�(����`K�쪍���j!�0�w8�q\�0�Sw��N;�$��0��ď���8
�������>��fਖ਼y�f�-�B�3e\��x:����Y9�H3iI�B
_Ujѵ��<�͈1ty,w`��7����}������'v��XJc �|�S�z�tK���� ����:�v;PeD3xu���,��۵�r���%���.����d�r��k�l'�K�����><�d;�M�W���6�����~4��N�=d���o{hw�!���Ny4�����9��C�[�]���u!h����sU�M�K?7��uDOu��m�[��LԚ4^3X��|�����7���[�����ߎ���13m�-GE~n�HM@�6��[h}H@=Ӷ<�=�0׶1��Y���N�����+H@�~�5/�l$
<e����>�atH�L�����X�<��lu�dC����	��Ⱦ���/a>�6`5���(��(K�/�`��U
<�Rw��*�E���Q����������_%I�ִ�
`�`����C�Z&P�2�5Ja^ΝO�S�h���^��h�Z�4�g���gsն �9y>}�K�QG?u����Q���i�B����<)Xl�ꌇ<��x��!����,�� �um��-�K�f�AT�N��fD����wi>�Y=��������=���cI��"O鰩��`)��ӟ")3c�6���/�Y�
%j��R�<�7���K$���r�1}�^��!cՃ�$[f�L��5�cL��^�W�s�D���n\l�)tz�3���SXG��ď����l�\%�=F �~K�>js"��������x�g�(���_�o�D�������~H�%`޿��v{̅�J^a���.����H��C.G�r>��b�U9�L�(�@��� �İ1����v��(ѡ��
f?;V��!�pe��`=�4=5��u�����cճ�`��_�vb�[�pb`z�F��)�j���3h���_���!kC��� �ܗ��o�KRj�����H���v��k����[7J��i�`�����\�H'_�?���qv�=厬��Iݍwi������E���Ll-���r��Q�3��*���t~�*�<���Xc%:ﮈ���؅�8Zb5�xRq'���f��+���a��"�<��m�"�g0ڞ�v�6�NI�e$=�[�E� �t��a*�:�(g{���"L� |� @<<�<ƉE��S�a����Q���s�s$����S�������)�@p�[$W~"�J�����h�yY��#� �﴾(��/*�_���;�zˣ�©�si�Wg�Ԭ�!����H����Ȧ�ԣ�𬶊k�d��l� C����Ɗ5�/�����h���#�#��s��M*����|�;b��4��P~|�i'��]n��G6��J�3��NCMA�J��:uK��f=�A����ѓ�f�}�+�4?��a@���X�M���?�]��Aj�\�n��q���Z�$ݶ�Kҷ@=���B�j92��P������w�e'1Q�WE����Z�Ë�ŭ�;��|���o�A�b"�c�6�z�.��V6�wݩ�$���%r����׺�^���Ta#�p����e��o-�7��G����u6jN�v�h�#�{��zEj���n���z����P�Q���)�����2Y��/牅=��(S��dxO|�#���܂����s�/��� '��I��f��NF)í��H�v�(�Е��<�G���Nţrx�\��|B�jpb���!: ���"��ʉI�#���J�����Oc�f=��8�إ�g��m����hǒ���\�OH`3��Z���]G�`毿�"��m�t�j������ ���q�x���]��l#�m��(�d��]S���r�����ԭdt	d�]������Sa7ۍ���Ӧ:�2�ՠL�4�Ӧ�2/�̛���4��ե���������+�-'���/GxH� �:����,Q���e�ZAj���ា��c�&��ZFB��&��$��D�[�t��/�O;..���Ϣ���M�]�f��eȩ�	��Aw#��ZD:�(��q �xM�@�%v��Og�2\����ݰ�Իr,�� ���������'��b���]���ݜʹ�63ϐ����c�����lj�0
�CR����'x���J���C�MA^w�0������Yp�a�od�F��6K�=��ٖ���LsN��ﭶꒆ���O����$�r��JE!��T�-�zn�H~���`���1��
H�{��4�.�Q�ȓ��B@�W��^L���/��/��t���_�1t�l���Y�@�f�*@9%-��e�kd/�Wn�{|�S�0���W)��A�	�Иf�-]JL�J:�ރh27�z���K�f��b!B���@�>e�?�|�-L�Gܑy˭1��8�P���'Oo3���p�CDc<2J���q��G�e����r��KQk�I]�'�LHc�2������95��]�p+��ܸzYA�9ᨹ
`{��6\v�s�˝�y
80��*�'�͒��}�����������}�#g5��j�r�-�=j�r(�j$�\�_�|-��@��	��5c��+ː��[��q�,��D"�����a���9*�B������Π�'R��v1}2�:VV�d�������q�xl^�KLLl�&�;|��o-ggT�H�MoJ�ػS7��/_��9Z��&����M���5���ex>�W��������ӽ��uE��J3)��
�@�G{����_c���-��`%n�b)�|=H�xtЍ�81�p�@�Y��^"хԞ$jL���h4�qC�kN�g�eo�P0n�jwT�}�9)��	4��I�}E�ڐ�57�莳+�W�Eп�$<�J@Z/]rRB��=B�������>ƻB���B��z��_���k+�3�N�M�n	v,�D��#�*5(�T1��?G�'pǲ/�( rr��&x�������)k>���jʛRޥms�����@��k�l�s33/�|猇���_�oaBd��8q���DE��,1��h|���ۋqzD���BX��#������*�8�q4�]#`|��c���������I_����F��H�����0��1�Y�
�,or�.����ǦFC����0dE��qn�0;�k����6=��f?4rs�O���'�V^��.��XV^�ւCJ�ИҊ�&~}|�{�g$[�̂�<�e�����G�c�e�X�P����!��[%�˓�꾦kk��&�b�M�m�߿q�ry�4�Y-K�r�-y��Y8[�sƙ�������/�5"N���`�ص2�����]����Cf� }%Ô&��NEN����y[,�cE�+���������+�2��_K�e�mٕLe����k��6�Zn`Q�v�G�r�Z�S�7͜��s� �ظ�ƝP`y�e`;)��ߡ�F��@uX@��]��kLi)l�@�\Qz<���q.eXL>�!G��iǗ���t���9�*=��2�A�f�*�nJ�:1Ճ��RI�xr�p�(3�7�JYD˵&�\^�'�o�b	���C$�2�3�Y7���q�l-~#���A�)�v�1d�O���s�r��	l*�پw�{荲����R��&:B_��E5�{o�E?L���^#��O�Ű���k�l�M��ڮ�A����Ӿk|��1��Ē�,���׉�i�A���>$��:���,0������^gR�����,���@���C^�%���U}��� �ȗ5B��013DU���p��6��P̮AfM[�m�� 6*�K5�M��@zxѾi�F�h�k6��4p�4�4�3�B=��G�Z���v������ZO���-�9����ҧ)���b�����n��y�F}�R&����e)�$�GJE���\r�2�������p�B���n��ܨ����2p�v�Jvy�Rޗe5�?@2W�f�F��ð������)�����g�̣�2��+�U$�u�*�\j�S�GzD*&;�o-�'?-���=g�4(���7|��^�R�?�'�pem��8<h:��	8�Y�w\�&�]�hR�C�)���X3|]�4�5�4��qG@X��[1WjO���`�D`ʒ܋KS��w�J��r&x~���ꟲȌR6�jIS�����q����'3���v�|����4��a\����G�,b���B���#ے2���R�$�q��+t,Lvx�\�Z�e��$!X'{]n�A�A�S_G���MAܦ�0²�����V��0f��76�յhG;�{1�u@���Z���!�s���6���:��ۣ\�[��?[_�A��5[�y�g� �JFQ����#��"}�g^wS�����x
|��)�%����$3j�.��H��%�䏈�!�b�����J����bqf�[u��,}�TP1���p��^Ʈ���L���x}a�<�fI��������2�o��K؄�O0��t�ߢ�8��Qs)��Y01}���w��F��fa�iX!�(/+rpWh���b�c�}ɴ��߭e@	J�3��`y��RcH��Q��^�㠄��J�n�� ~UC���t�j����P o�2��V����Q��u)�=k��ʾ�����:�䖦��ع��
W o)�	�L����U�'t,�X�}��Ӡ(���7��{t��Tij͡��7�wyz���ԔY2;2�︛" pbECٱqTAw�� ���Vp���ACun�eji���š��3���@;�m�:�"=����l�cn�Hű��e&6$��ɒ�?țn�G���b��3�c� ��iD���8�.M�/� �, &��ɗ���7����	�F$Č�t\� 9B>���$ ʁ~��C]Ho�j��4��ݶn��m��4w�-� �$�>%e���<�x�4���3Tm�YDw��~^#���c[%��D���wҖrj]��.2���Ϲ-r�����pIv�<�":R��9��ss��yQ��3I
ر�nn�����|������0V�u����Ɔk֬2UT��pi��p�P;��*��%�j�'KA5�=��{���4{��vƂ 9���z`Iw����N�5K�jL�jϣ
`�kA5�����s�ORPL�c �Ö�w��ҔB��Xb�Bk�\���m��?�&������5�Nl?Cgؽ+ ��x�~�]������8ԟĒoLf4��\�����0i]/���C��2���nd:�ˀ��3���9u��	�/�� ��ԁ��l�p�����W���~!o�X%�&�C��s���ۙn0�B���JӼ��c�k&�z�6Ծ��#��B"��J���|.���5D��'�;��"ڇ�ݰy�m����"�ß����Ţ��nvn)aiR�L�L�N�m�c��LpB@��c��C�'��I�av$���!��#-8�BF���� ]&�����MQ�Rc��7"����~�Lk�!{m�k�i@N4UM^�l�KQ���$ۅ�Ou��bi%*B��(<���D���1�B�hX�V>�;�'1%���$w�\nGM/l���{��A�ߒN  >�RՓI���Y�RWl��%T/&�jà�C�sS�����"�	������+v�,�
 9��.�o݀ۦ�ڮ�Ɂ�J/����O�o�
3Z�u����U�T�-~�$7\��Yߝ:�	m�x���J�oF�nx�o���&�w�N~��_m������e�c���	fՃd�WY%�Q�|o�/��`7]r-iT��m����j_D~L@���M"���V%p��{$��XR��eu�'"��:�b�����o�?�W�='f܎o�n�+�p�O�Ğ��
�("���]c�7�
�(�B�Y~����[}�H{2���x���0��l�����9��엱�����M��_4wt���ޓ�X:�$n|{��#z��9����9�&��)��M�7�Eet�#�]�����ޠ	��_�:�)A]\�X%��Z�I䧨���ԅ�]�v���(����xZc٠�tע���$7tZ"������Я����e��]ͥ��G�Co5,�l��kѵ��F�A�(�"o�WJ����#�3�NRuO��\魌A�۰fS0'��o8ᅱ�mh`y�a�LS�Ҕ�����?��ȿ �CϠ㭕$v:�@��'܍�k��S�J.�p"8zw�1O�I�N�3�Q����5!�,!R5�nU;�&
���s�c ���x�n���� ��e>v��Y��"�[�Q���z[&C�A�i����`�����)��A�	�TJwS\~��$��~5Y5���&��&j�̌�
����oT o9f���7�N@y'"�����0�|T�Ԯҧ�p]K��|Nt���Sn��i�[�H�G���`ٰ�$g���{�Fu9�¨���(<1u%|!���z~��l�b;~SJA��9^�#��v�b���素�O�],)N]�!�W��x�pk������g��<1���9�O�~@`����oF˯��s8��H$wXn���{F�6Z�NsH��gh*��-���=��/��X���,����r��Ŷ�rf
���Tg���q�qm��]n�;�.|j׋��ULP�M��,1=|BA�<�s����v�#L(�%҄`)
�9#,��q'Q�=,�}�ws�Zb���!�t!��G4@�ܦ_��o�?~���*�3�(R�&��J��%��dC�q�$�;���	r�E]n�[T%!���E:���K�:���T$�	�{����Ԗg+���?'�{Ɋ�?�R��� �Yă�o/���)�D_�q��=�c�9�u�hp���K%�'0u.�C�!c�#����5��c|�qͻ��XqS�O��"M���7[�h�O!������asVvW�6o�l��������B٦�]��0���}Q?�8�ibjN�u���/�F�i�kR �qLm�67꒮�
4�}ʭ���c?c�S�\��o��/.�%��h��)�dj��YS�v͸�;
������_��
,z5�B�����|�+Y�����yQ~J�oU].*��肍��x$��T)� �o`<��W(��/H9t��TCjŅ�,%&�@4�x��uO�U}r�0�QA��{|���nH�O�	�ξ��"���%�h����S�;���p=�`���`!�0��&=Q)q�(�'�h����[�*{�����O�-�kA����.�R���q����6���.�!;���V$�M�>F�ޘo.���)v;��e l����Tp?���