��Y0SY�SSYP��Y+SYYSSYQ��Y/SY�SSYR��Y,SY�SSYS��Y-SY+SSYT��YNSY�SSYU��Y'SY�SSYV��Y(SYSSYW��Y)SY6SSYX��Y*SY�SSYY��Y$SYESSYZ��Y%SYFSSY[��Y&SYCSSY\��Y2SYXSSY]��Y7SY�SSY^��Y5SY�SSY_��Y3SYNSSY`��Y4SY�SSYa��Y6SY^SSYb��YCSY�SSYc��Y9SY�SSYd��Y:SY�SSYe��Y<SY�SSYf��Y;SY�SSYg��Y?SY�SSYh��Y>SY.SSYi��Y=SY-SSYj��YESYnSSYk��YDSY�SSYl��Y�SYtSSYm��Y�SYxSSYn��Y�SY=SSYo��Y�SY�SSYp��Y�SY
�SSYq��Y�SYSSYr��Y�SY
�SSYs��Y�SYSSYt��Y�SY�SSYu��Y�SY7SSYv��Y�SY�SSYw��Y�SY�SSYx��Y�SY
SSYy��Y�SY(SSYz��Y�SY�SSY{��Y�SY�SSY|��Y�SY�SSY}��Y�SY�SSY~��Y�SY3SSY��Y�SY8SSY���Y�SYOSSY���Y�SY�SSY���Y�SY�SSY���Y�SYeSSY���Y�SY�SSY���Y�SYtSSY���Y�SY�SSY���Y�SY�SSY���Y�SY��YW��SSY���Y�SY`SSY���YMSY?SSY���YrSY�SSY���YtSY�SSY���YsSY�SSY���YuSYSSY���YqSY{SSY���Y�SYxSSY���Y�SY�SSY���Y�SY
�SSY���Y�SY�SSY���Y�SY
�SSY���Y�SY�SSY���Y�SY
�SSY���Y�SYUSSY���Y�SY
�SSY���Y�SY�SSY���Y�SY
�SSY���Y�SY�SSY�