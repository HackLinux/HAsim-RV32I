�fu�`�t����s����u$2'����c�ID��Ƃf:R�T�,��Dp�r��R@�yIN��o"R��<�
�r���|I,ݿ�an�~4"5u�׃[ܜz��]� r�h��X7w�%\Q&�'lk`�����0)�[�0d���(�lA�K��,=&A�Xl�Gl���L.iBl~W�q�\� ����*ʽ�x�^n��	�)���p�=Pdm�}�&�Ի��6.ۉ�����+��H2"ԅ=��t-F�\:jC�~�u���S�]k��3��.�3r	B�3�T�YL�_Py%S���L��(��xU�^���y�dh�J޷�$��������,6�j�z��[�]G���e�c�m�k����Ӯ�Ю�xJ�ɨW���^֯˳F}�����f������*a}=-*��U�d�`�;&��g�����]����9t��/���w]�T�����J����%�ʳT�S���ƎK2"����Y��Y��;�+p[�>�:	�,����7!�n4;�5d_�O����Lz�Z��P���5mvţcn�Z�B��V|פ��ne��,OjtVbI<*�8�)��Q�uBY�uJ�u�K��69�xґZy��Na�����<(>w#Z�)O�va�P�u�҇i5�f��?��FmTy7�KUO����n��S�BWC�8��1_�5_��.y<�������rMe#��")���Uc,db�����(��f/м��&����6N�����^�;W�f�������u-��5X�(�ҷɝt�Ø�`:bАL��y4��Hy�e�	����IЌ�%��*V��W3JRa�9��q�V��:u��虴n�7E��f@`�r���Q䩠��m��2��bC$�m�:A�I�����|�
�[Q~�:b�tpz֭F���l[��f2��J��K����Jx�-E����c?g*�60��G["���D�(9��O>�l�
�����Ʀ^&�|�d��o+��i M��q�<��פŨ�(O��c�'_x�q������q��><ת�wA�����ʛ�eQ�=+�7*�<lN��B?��VI~b����&=�k��$�&AJe�"���p��Fc��I>����"zB�(�x�[�BrL�-�x�Ϧ �lI9���t4�8���Q����餩NIS�cj��7=aԪVH�2	�oհ�HkxM�D5W���ן"z\���Q�4�A��cV�|��x��y�+�hm���SJ�#^�;%��"3i������`��/f ī7('��o��Q2p���B��6ӌ��I3_Ҥ)��}��(�M���p�����rNΗr6�晽r�<Ӊ���^�;z���z�P�V�=��Y!��A�gGA�����m_7������SnoeY����Z�3������H��,��vbb�
��k촉uć,U8��:w�Af����� ��̋e��C��������y'x���ͼ�b�̛�Vځ�T�m͕_<�6�Giױ�eE��9�D@��ض�Z�畠/���T���`�I��r���ȧ��;���I����I6xҌeA�<.j�#�-D��:k�5b���Ҙbt�wm�X�+{ue�-<8�ֵ	�׏=q�c����+�kӠ4����X~h�����DE��*����#�OjN٣6�@J�]M���������i�G[Hܙ�0���ҕ��h��%6[p����xfI|G�Rna�O��x ǎ��]���>��2O����\�(��_2w04CXE��/wd޷ t؜<W��^��Z��[�(F1�#�,���̽H
�����
��`�훸7��u=���YF������`]���	Va�OA��$4�aq����jR��棙�qJ��LF0�^�Ɏ���j"�JB7���Z�?V�H%�P�T�zr}�1'Pp��bx�%�'+Q�.4�=�t�m����[��b�eq�6Y9a�^1�l����:H�-�.ښͦ�RΤ��E���MO�:����!�1�B�UJ}@3p�����J��J	�<�F�n��`&5&K�|'���[��^>�&T�T3
�!�_�ԹsQg�j�6��ܹ<;W~�����S�s%�����8��U��N�iʚϜXs"�Pu�Q�v��v��S�����Ā�X���"�Xrޙ.w>^������&�]��L��I��е�tD<�@��@}E��
��o$*�;����(I��@5�C��֎a�_�Y	V~�!2dG�b<�Nڭ>d�V	�x�x���Q�Y"�YI���PL�c�B�&n��b�3���]�m�CKA��� W��������RV�zYF��ǻ�	�~,�q��O�	�gN�!�A���C�h+j��:�Y4���*0R�SU���IԽQ�b1F��j���wB'�����Mvfԭ��p�v�n�ޚ�`aͳV,�����D�� d }$^��wXy{U�"NЫg� ���O��B���;�]��d�aL!96����6V�>�Ӣ�ݕ�pg
%�h��x�k;�:�)I�����:��[�H� ��aÞ;'lgݒi�`�y��2\*9ur�Y�N�m,6ٽr)�Jt�f�������3�[�k��4����tB�#c%�4ӻ��ق`b����x����u�W�XE������p�J�b�S��3cO&$4�QǤ~�R����V�n�=�0� ���'��%��-�h�SjDr�;���.�v̀E-6z�H��oz��q�Rqz�^=�_�G�q�r��`�����k��-�u�P� r���g6���eo����<e����~�+7��K�~Lep.���*f�K�6i���+�)jF��%�EM�(I&/�M���HK4��nf�[���+��Z2,���ښ��KC�}0����;sZֲ&6P�%�E��lm,'�l}q����%��ܰw��kڟ������/V��'f2��_;M��:U������G��N�/���Π��Y�X���{��L�3C�p�hd�y��)�V���]�؎ ͚F��������@U�l�)7[~T'�|��=F����=k��)�	��|�:GS��E��˼\��ZŇ�Y~m�ǩi��kc;"�P0�%&%#�#M�k��#���$.Aʹ���F���0�u/G�@W�������)Ty��#k�J+m��H�f�J�����?F��4*�:�s|���󂤗+�	�<x��N�N����g���龪��|�~q�+֧���A�(��m�L 00���NqP�ؔ�k�d���(!�����t�q�pN�,A݄#+QY"tu
wS3����M�&B���#��!��s����Q+����G)��^��Ҋ�"��G��]��3*)m��g(g{��>�Dw:S�Ϩ{J�Ԟ��/u�n@q���h�V��q�_�8�d���˷�|B	�{MK�����zhU�Oo�j��)����0�b�?������Ӈzڐh����e+b��t�5_Y�ϭM���������Pō�9�?鳻`���I�p�=G����L������ k!wޛu<��e�T�:en��%8����)�Lٗ���D��Y����"s�[�"c���)~�o+Q���綛X�P��߆�E���}��*1#T���<�OI�V�qn平R�{��q�c�"S�!���d-���͆�h��x���ζp�u�|t�-[�_�sʠ�kKI����`I
�n�c\Y���hkp��	�ά8����1�zˆ�G�o=;f%�s)C����,��x>:���2�GUT*�Y�F*�ڳ��gg��^a��<aad[$3�ɦb(�~X�f类�����n�k�j�la��.N�SrW�h���)B��M]�:s�;+���_�������Lb����:s�:���NG������#3w�w����l��w���R�`��mh9�Ĭ�*�D����m8~��8��P"�$@;S(6fqv�v�hd��y��[,��s�������U�'�i��j���=�m���3]XQ ۞_6�3(�1����V���:BKpP��v�!w� ML�^�c�uUM�e&�Di�_��Y�	�A.b03��͡O�}
XWz�@N��K��\��8��F���.ĤN+9���s�D�~/��t�8��SʒlN*�0���˾�'�ÿ�̅� ܁�em�AfeM1�	�[�o����Q��_�	����-2~� ��e=5�Y尝O	�g��m�jE���ᑇy��9]���:�:�al��B�+uv�,��#
c�c�M@�*�9�k	��>��Mhw��
(�Wg#�ǯכ�-.�,�]��<Q�&�������sY�f��ɛ�����~4{��������4���l�љ�z\���s ��O]+ �T��H���t�ˍѵք���9����Zw�z����o�XLɋ���N�ؙR�L��=lP��w�.�  ����~>5"�ʝJ�I�3�˝>����\ɢ��n�џ���P�����s��u`P_ �TN89�pAj���7Kp�ʟ�^w�o���;w�Ъz��H������,��k�ˑ��|a��W&����e�@�;�\�)��Z��A������n���
%�xX�J�W-K�`�W��%�?#RB�ޑS��ֱ/�o���K% �u�,6��F/ur���*E�]uﳧ���&�V���Eĺ������L�h�Kϝ�w	�J����L����*�W�J�a<
�D,1��5�5M�'E���;��Ǡ��.8\&ݻ@����7W/Җ�kV�|���R|u>5ŷNM]��LY�=�R�5C�{��_&ZU�2!9@�:��S.`���B�1���3|.�-E�����m�^1~�D4�զ�����&��Vᵡo�_�5��k���U! ύխ礦���
g^
.���� *J��5����Y���l�*EX$l|ywČ&$�b�)��3���C��
�������^����OTh^�x��ZT����?jT;�v����x�*�;3q54Bp!�Ģ�f�$���o����W�4�z!����<N�N�f�.�-)�u��to[�ٽ������)o��Hv�#{��Lq�fMI�_��d�	����$����깅Ø6:L�HU�v|�֛��#���|�Q�)n�G<3���g^P�;����̘!j�)B$ �gCv<�}��Ճc�J�g ^D�H�o���Al$�6:�*�y=)���-�/zzvZ��nxj�b*�����k��ԙ]�,�9V�] ��T�)*G.3�Z���GkQ�3]z}܄Ӊz��>���1ۭZ���?�y�+��з?��[����`��M����P�v᝜]8��eߊʉz 7����Q����0٦��gV�v�J&,�3s�i�	g�I����'a�O��B����y}��5�;�mԮ.�&	��^�����d:wqkƛ��k�W��+�y�i
R�z%8*f��D�ߥ�s^C��^��ݵ*ƴ&*�uږ���#�f�#�m���ZL���.�k�b���~'�)q�F���D8���~>SmXڡ�T�֓�L��lV,̅Kƭ^.N���f��]Ԕ���ؽO����Wm���2��.i���T����,�x��+��1��l;uf��<7B�����EϞ��Q��ܯ�a�R9�k�3���3��U{�j�*;����H���C^����z�d������D��]OO{��WȎeA��M�(q((�G�c[�%]]�dF��"�R
(y��5�@+参O��v�tdp�Z�Б�Ȁ���T�[�UF��e�vQ��	*�֕��%!
���L��0׌����Z� Ŗ�\+�I���ۋ(}����e�J��i��2M����3��i(.�D�c�O��Z����{QӸ\кU"���	�v/���^�E*�\�QܾnZzѷ3����>�
���J������g�
i�WǄ&��
���^��J�6ް�J4g��aXB��M���3���~�,�P�n�B��G�g��W����&Y�G��o��v��;�E���_��	x
�D�2�j�,��̀&F1#}��)~J����(8���߀H���lc�kdb�k�|�Q@�o�|x�;h�mA�Mi��m�0�6{�n�
#�fN�Fp[�d77d2��%+�����^��Al.��ӜKp��Bp�V�%z;	: hd�3(p�������l|(����;��m���|^�`*�`J)�<Σ�{�p��� � �dk��KW<�*��@<��>Tj4J�}[���zO�?�:~K�?�Ao�u�s�V���$�rK��x����~�`0o/([޿xA=� �����j��/p~�����:$�t����`������.;�:4��H�� #��L���!�-�TNs����C2\�^����l��lS����
�N��o��/���9��?g���wy�}�i��fqZ��j��#p% �J�h�M�,�'�0`i�Vٟ��z0p���qU쭭��JN!���n�U�I�=�Vi_3 	�م˞?V�T�}6j�?h7�g�\� ���+���Pq(,�f5]$
?'��/+[���z��G�[���Uu�̸Uyb�q�e��.z���}���к��C۟�}.�VW23���9�č����H�q�0"�_���o�a�/��N��S\�PVΞ����,��5y-���X3Q��D)"o��Y訖�	ň���1K<r��ƌN�'o�F��,�P�,ԋ3O��� p6,m��^� k�$��[�9:tl���x�6��%�UZu8EB0�:�k����qJx�)� ��)@B��	�Œ�y�Yp 3.�!�M>�:�/w~dT��� �%�֭f<ܻI��B��;�:ڸ�.�+JV)2��+����#C�E�(�f��q�ÁM\�w?���H� ���v8�n��i�qF�F$�)��Ά��2fq�� p�L�r-K�iW�f�E�=�C����*h�������g1�h������.��n������.��.���|lC>�0V���.Gbd�s�\����}1���H[�&�Z�mu�XQA� �ޣ��e�մ���E��v&sK�N�	���qP�P?q�g��+��{=]J�'�����>�ՍF������U��\�%����KWČ �9w�Q��_���炀������iݠ����u9�� ��d�~o��F&�7�hbq�A��;��Úu�]��e>,��s�gӛ�5�Ux�gEiF��Vgi!Մ��y�a�i��4�L�'N��_�3.Y`:��!�HgP٬�Kp诛�s�]hB�������'��+C��S��LRW.I�0v��2��%�}$����PbT��i8ܴP�u��:eG�_�8/x�4mM�pϴ��"7w�S�yH�B{3R-� X��9�콽�=���EX���(�
����e-��˨�1Ļ��ae�0�|2]��jK��:�S-�g�e���u-Wv����E�����]w#{{w|='V���q׉�:^���7Q����5M��,��!����R��Y}����6~�{��C�Zl��_S��՚�����R�������2v�E9��e
��������y���t��C�&ø�j��c�t+����V�S�:����s�-ǇTv幔��8��w ��o��OԾ�>X��P��g5jN=��eP��i�R[�dZ�`�+��p�����}��c���p���-�VO�J�e��e��T{k� ɞ�߲nY양9{eSx���l��r_��;	S� y2 ������(��(+���P��IU$�<Pu]9S���Z��s8�h�����#E�����S(�g\Cx	r��+4���P���`�[s��c�P����+�D�cң����jz�V���c�fc��х{��_q�B��1/�ܡZu�C�䑧F��x�����F(@}���Sä�����}�:mӂ��\</rT���0η˧����i4zf]��xC�c��Mm>��S��f�����wc�j�`څ�_���Q�ST)ry���uNi��y��Sgx�N'm2-[�8���I�_Yi�z⼻gRZ��P��\�e �.��)S�c���.��+�]���_�M������@
�J��j��zċ%$w�	��Y25]>�Ɍ��� �҂��OM#Om�w�+�s����wRh��˯:���TM6ѼC�z�{�w�`C/<N���*�=�,^i��H���S���}�fp���wO,ilt�S��rt��L�ᴇ=>�F�=��G���\<~䲇\q3CAy%�p��-���St��E�4���tv�X�҂�����ެ�= x"����h"��o��3�fD�#��%�)�c1������ta�.}N�Z�������C�@�z"��i6 �f�xp�������-�[I�'�*ڀᯰj�%KFaBC�Ҷ)��Q�nv��=�Z�����qj����SM��	�oT�ݓ]�+ji34��������K�i�#Iy�W��|���۬an��T/}#4���{�]X�7�^<:�2ܸ��&�=�/�#�o.h�V&��^.���GC�MD��������{��[O�\Do$�zƥ�
y��kW�Z1)�q+��u�J�kq<���1���(N1+�S��ּ��-z����IT��#���*�s����ęqj�r�f_��=~]ܿ�]�qf�UY4����OM�8k���C���x�Eʤ&DфZ��~���H�c�J��q�_���	.��k��<� C[0"��Ufs�KJ��@�h1����+�G��I�/�w��M�V�Asvx��|=b�O�]@J�~٭ԙ$����O6 XJ�;�Y��ՙ�M&Щ8M��nj�j���*����Z,�Z5!�5�DK޿��ܵB�pK��0�Z����C�Cz��Hß���8;	�N����D��8�͸\:$1�F��������Щ��K�L�Ulv�����H������(���{�%k�p�����^k�ȏ2��?L���hE����{�=7J��C%�܂J���O�bo�����'�9n|�����@uV��Ö'�̰�T;)"x��%�z��)>ړD�]p�/~���ݭ�v�a�;���չ/=���w��^�n��*1�S��aR+5���;w�G�L��\Dp��L$�$�\<a�3r�Y\��J��	+��/T�S�p���֯3b�9���*��E�RY��5����P�k�Dܴ��	{#t�^����m�19EE��L4<K��\g�T�]�}��6����u��}���x��]������|,�sS�,�ZyJ�3%~��el=��h�m�0�d����^w�׆5`r��Uh�R� be�'��%��k�Ff4��roM�b�� �[d�/�l�˩A�V.�>U+�T+g�yM�a0���U��V�=�&̮^���+�	6!�T��p�ةSkGR�1;�,