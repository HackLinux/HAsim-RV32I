JٮCH���߷[W#��B�����}L\��)Z�I P�,�06Y0�y��e�%���f���� M报�B3�rd�3�c\���)�e�k*�$�0ّt���aj�r=
�k������2ҕ�^y���K�u]�]��bؼI����:��_5����lr���X��"��m�BW�l�� �荿�k-�٧[ޮ������xb|�,g�d&4�ƒ�|�W{h9�j�� UM����˩��ǵ�����
�v�,̢�W�o��r���g|��5&5I��墮�_Bꤧ��q��NQ��1�}�̅�|�BS� ��^Ն��DzF���5�}���[}V���{j=�М��pE�v$m�g��~9B~��|��z���x�Ԩ���8Se8��Qb�?��J[ɰ֭��i�a1�:��cU�,��6���1��	[�G]�/�!SzU�^N�U�DQ�'���;�
� �	�J�������%���ANDsz�O���HY����sfv_]�D�׆h��9�Ey��[��˖Xo��T���U+}�,���(�K��t��"[�Q�;a��7Cy�̥3qq�$�7F�(b&� (5��$E��E��7��@�l(^�Y�@x ������i�5��������x�Q�@n���Tf�	Sh%J�+)u�oYn1�nw�P�|ʚ._��1z6iY��IÀ��e�m���c��LN������d�X��E}YΠ*�\�6�r�A���$3'�9����ev�i��=�T:b@��PG�M���lb�ɔꩁow	X�h���;�բ!�^��otB�N�'����_z�v�u
$���V�����d���;�'���y����a\�0�#�e���C,2�|�Q&96Z�{2656�wJ��M/�`�oB��*��b��T��>Y��q��YN�7^>E(%7L72�����n�S�;�N��G���t�%�'����m��o<^YG�Nk��z�(���P���&��ώ�� XL[Xǥ�E/���Kozj�E����MOD���>���dT��?��?�q���>�V ���0��#�4n	����]�<�ɍ}���[eJ�P��Ch<�g7��qdm˝�e�̓��>4{n1�Vv�S�e`,H��:/��~4/��%a�r�b��u��<<�6pl�iy��E4��6��9��Z���T�cJ��|V�-��1�΀��j�b�2���Q�g�`�SC���\�+ �o��k� �T`�Bd^3�}��Lܜh��~C�uPo���G-@j�S˜��✕	�/#hE�v_چ�����m���Y~׹��[�^�T��x)z�h|���cL���L?Sq�S��!�y|�Q:���"��yaOǅ;0�*���:<E<��� ұ�!^����v�i��'�����-U'8��۰�����Ѐ�jKZ<D �@��,��,�E�oFևM�-���6���d��|������ߘ���ҿ�@�[D�$��Y��F�����c\�]���9���_>|@��SD�t�2���W��|3�j4g�m'{��]-�ɧ(�8ԍƲԀ���J�N�s��3B_U��©�KR�͞��1�O�"���w���<��b(=�h��Đ�p�W}�'����[C?���Ϣ��G&*�H�1U�p<j�ޠ,Fg��֡�h��S=sߩU���r����\���܊b��3n�6
0���,��i�{w!˯Y���?=����x@Y#�d���i�%��췊�x���F�X�`���IC0	4� ��+���_"��@������X�G�#(��H���$3�����~a#��}�[�g������n���u����W�|��9UE����A��*�z~�| /pS�QPX�2 tL6k`O���/����$�N3�=�c|	�r<���I����h;ERMqI��6M�w�Cw�Kc�z湋��`K���v��)T²���V�o��-Š�m��[bDjt!��ڰ�`^Τ�`S��
Y#(�𷮎ޮ�_x,:R$#L��'OվkJþB f����`P{���Jx��<�Ϯ��g�%r��!��w�`�c}���,&�W*��X1t�Iұ�W+}��3���bø����	�e���(D���
���*�9ԯA����~���}�.b�	��;����ep�tZsL��>vw9�$��E͆�zM�a�Ȗ[���L����^l�f�n��<�����K��x�o�D_�K�Џ�_���`�.��NOP�� �!��%���E!К�n=��y�G�j~]Q)3�����F�y݅��ǲc�I�>��~��8�>V�8�~�Ry2���/��ɾؕ�H�>s���s����L��W%�o���,}�3��ʫO�K ��3�TKHh�����&y����?N3K����z���kcM��Xuh.|z��Uk�q�j���A�ɔ��i�q�Q�|H�ǅ��zN9�S�wfa�e�����lό�}�^�`	#��6�쵆���M��m����[Ͽ�FCq��B�Yi,y�>y����3����4!�� ��°P�D��ک}��-�c$�CN6���;�c� n����= �U�6����zïn*fO�	�`���F�7"��*,v�dd[�ffo�F����������{��0D�7����f�w3����X��G��*H���kM�~JX�^R7i���y2F��A�[��Anݐ�:\��j"��%�ֱH�,�kgG��[Ė��b�������7v�2 |	����=��#�(z�{��o�����c��<m���$*�iӔ���k�-ŮJɴ6�%�8�4�m��
ENE,l=�y�^Z9Wp7�n<SC�H�oD���/�D��V�wh��zT���6e_��+p�E�@�ʮW�K������d,�f:�y����`~+x��7<��{��u�y�=����(ނ}��/C�:/a>^��ܳ��籌���N�UM�19���`kB�&Ba9���$<��HX`9['�%�d��[��k����^ʜUR(�Q���Mga�xZ�i8�#����b��e��U�킣����}u��s�ru4_�h{Iyl�1�[�}q��.��/�5a,�t2һW�o �&_V?}nw�|�<�[<��
z���7�I~����S��F��r%c�����}|Y96'�����1^m���!��)SL"`Ca��E�U��Ə�[��'��JC:�V�l�D�?�K53Ҫf��UZ�^���8�fCյ�1�� &buV��\Q	�v��fz�������1���c �)��9� <>��ud�k����N�RU���|�Qk��(�r�A����y|���y]¾:R�k�ug����H�?%���(�e�t����z�R�Q����@0�O]�?D�Υ�,Y� �2L~!������f�_�Ʒ���9sș�̿ͣ_�9�G"�_�e�$X
�B�l�c�<%��\�u��_ݚ�kk[Ws���K�SD��B'M��"�|�4j5Ql�K��Yf\Ete/�gn(b:��"�yL��(J�
����|5Z����X&�O�c�0��2�'���`�C��8�H.�3�y-���;,�7�]:�ֿ������y�-��!�<H�V��n��He�f����';+��u��)͚�tm��N�Jf�`A�6�ҥ���W����0���W��k��60N�
Q3�Xj�+9p�]�f��!D r~�S�л��"�����`���y9"<��,�$sSU,-�Hf�f:�F�����)T�E�%�ix�R1x� 5��$���. C�h�*#�̝d)��*T+䟃�;��/���t�M]Z�q3$�u滥����Qf,�h!�_��ֆ����/V��~��%��h:�H�少SA�%p�b����;�|�{����31!̞���YQ0?y�_�H790��P��[��˳3c�]t{�]v���3�#]+zN�p�ҏ��{�{tі����A��H�ǉ�g,4�bD��ф�2�(@��w[�-e�������W�BⒼ ~����?z���
?M���O���,�+�����hDN�>��si��N���(��pc ���~� CQ�k���8�66��C�I>�{�AӺ�����u���ྡSU��m���%�z_Úl���Z�.�h�9)���.�������+>}:X:�	E$��Z�o�B�&��#/(�* ��� Sʤ��Z�,/&��|z�t�yi�����'O�X��L����\��̍Cr�r�&Gs�yR��-aR��+�a���@��$�S�W	����B�c�~��@���	?����