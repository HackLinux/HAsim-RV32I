�����;O�t$ jy��s�����X�؁3�v�E'�5:4Ģs>^Cg���ű������O�~[�`j��Jg�PmQ�u_f�'M�y�4GC�n��×��YʰF~�rq�zP�&&ڙ����[����sп����.���+��}ˊ��p�Ixwi�1Č\�f��L�W���b��C=8߇G_�gTt]�Ǎ�j�CVһ��R)�N#���oxiF^4a�FV��ܣ�L��#�ˮQ ̊�;6qC�"-Rh�#L8n�7�e���k��<���y<��z��<N�<P*֊	���΢5�fќF�&��	GL�*щ��gI��/˪Ld8qm�6�y�i�q��1�Ӵ�Ckh�v����p�8�r���qN������rɏ�k�\�Fm�|��K�v�g�oY�-b�Jʕ9!g�s�ɱ�4�uW^7ʗ��]��
=����I���pV��@��EO��ů�Twv��z�Ӟ��m J���Rum3'hm�9R�94�"�nM}/n\��DG)��=	�%�[���E[E���c�c����"'�2<Y[|N١�F[~�ߝ�ąE�DМwp���`�"7Fk���wٗ���d�%(&2���J$�`4�I�1��Sa"F �"!�!����(��)1�IC�	2�ٔ���bi M60͔X͈ɦ���Rca2h���h�!�d1 &ʋl���RmcQ�JBQ����&fQE�IDkdC(1$���Q����Ěɢ�+�J�1�ȱ����k�KbŋPTlmF��ZBd0�Ѣ�X�E���h0EKETkF�QZ��E�Œ&T�Y6�I�Ƣ-��m&�mk%�lI�Tm�-���h�ƨ�$֍���EQ�F�[E�6�mF+EV-2�(�5�5�EQ�Tm�-��Y+TTTQT��DF ��E-kj���Q��,��1%�$��#QBa#ģT�ƒI��-d���6M���!06(�4�0�b�37�[�Qc
�G����_UQ/��To��>���˝i��j%N=�q*ڌ�9BU�+��z_}� ����);3�$���\B�����f>4�ۨ�"�R%N���Em�����5��S������)MAƔU[T�k���g	)���?����z_6uG�U��z�����L�G)�n�x�cف�7��{h+������S�eKTq���.eht���@�ix;��? �z:v�*(�_E�|�eJ��SmC7f2c��;��=�LK͢��ע��fZ}��6��h�s���8sI��N3���߶������y�O��W�;D��E�/�k�X`ow��Vhh��~��A�����9A��?YPbOo:9)Q�׳R}�3�i��jb�|��;=c92�C+��3L������Qjε���B���TSLm�T��n-���]]Z���o