��u�U�.q�~{i��~��d���&=����e�խ�O^dH����C����B��� 5�̣��󯇁��� ��@��/@�q�+����G{ �Tm��mH��-n�|�?MG^�/�5�ۇfP�O�G��dc
3�OnW�@;�b�����rEPA~M�cÃ,�|����q噔cF'����(�$Ҡd���p�>�I��^�e���=_�����ZѾ���\(@���6 ��9��G���9}�a�i�0�ݸ33Q�ha���v���R8"y�%_J@E3#Hq(�J%��Zڕ�[y�{dd���T=E�=�05"�-)T �<A�h|QÜ�1�=Xx���H3��D��X��b{b���T�ZKd[��Ǚ�/���ёX�KU��0�Q\�
�r,���D��ұc5��өa&�'Szn1�����]�7/[N"�/g�HN���)?��������i�
j8Ģ���Hۋ�nE�;x2s[���v�j��'7"�A��6qw��&7�{���=������y����EG�2�(L�8pſ��sA�u-e������X�/o����j�$�$�(��Qѐ��A�Ͷ�qp��䏘�=Ŋ����(��n��8��W.��9���-���
䣋��^���_�8��;S�T�(���"/�Pd��p�X�5��N�9�k�Њ�8R���=l!��jے�*��ȝ����OJP�`�%XN>�+��7Y�� �3����B�F	�YJ��65���Z���k=��I:����f�e}�c�W��?;]�q3;�Z��pO<ǔW������PI�gP����CpSێ+A���Uk�m�b�|�w �s��^���_�ہÜS�4sI�����[y�a'���`8���K�x)�2M�y]��*�E��ۨh��#G����̾q����EJ��螵q��I���E���(a�r�WW���m hr0�ikU��Oe5���Ǌ>���S����Ӡ��#����i�6�gs��L�w��ruUz[3�V)_���wt��s��ڊ�5%1��հ�S>B[4�HQ?��@ќ���/\�	��ڏ��}$�p�?$�{7*^����R��*�/!�K�7�U�u*T�Jx%*x1��7��Ω���6�8&�(e����纭%�~H��?���T$�v���
Һy�\�k��^������7�ǽ�+��fEaT��3T"W��L��8�<�uEny��ᦠ��0e��ƣ׹ P��Wp�?��T����Z�?�m�ò�v�ֽMQ�?�� U]���݆�����(�5��~R.�0������f����탛�'*=� )�F��Q��,̭�@��-�삨.;�N.���Li�Lkw �78�>�<�G4��i0F�Fk�?Ԁ��\�:8x(-����_�Nm�?�p{�׀�3:
)�|���;���N�:H>��p�ה�r�^pW|O
��=�5���ŋʊP�%V�͍ԙ�9=��
��i�*�Ǐ/����HUЕ��1=�$��;��ts��\�0��Ǭnm����l���D�=�����QS��3�p�V J�w��Ww���2�W���]�C�����/[�N}���sw�l�����R�S߂�w��] ,f��.����g���b��OG�x�`K:�?���>/�3YOwt���py�����짝�g9���Gs:�1A3��Тz>��ӹ��gvR��9�s�i&�}������'��E�o�Vg����n���L���z���N3��Rz\ik"��f�b�Ǚ�����띕�4�ws�.d�����oh;�g0��x�����E��e���Lk�u-�U�,�ݞHϽ_��>�
�=+���u|v �:�l�r/%�Wi����ٱ�Յ���9�3����������Q��+��dC�@�,�R0���qC̫�gK�{�U��%��u��@��L�V�j��$�$��hj�q ;��('��P|�4^�`+��9��q� @LWŌa���)��l��_ �#H�I�)�Kƌy�K����m������g���;���c�����}��u��?臣���^ԣ����>�#���9�	UW�qV�O+���a�M�$�F���-��1C���qy�@H�$˼�*�\q2߿����k�IV?����]�|���6TE��T����sQ�����=�Ǫ\cMoO�R[�#��{�W��1߸�ü�TXe+Wr3/�^q��A�s����'+J��HpV����s��}���d�q
�xzC��;�[�іp�?cc��iu_�|��[�2�����N�n�\�CTS[� 4���f]����I�sf�g�dbNU��:W�����2�b�F�. T�2!�qF�hu��nTZu�`(CO�EBs\"���b��Y)M��.�3dm���Lgq:��;�,h�f�������{ݾ���{���y�DG���EE����v�����z���OF�廎�㻆��Ύ�����of�<�������S$'^R��>�2q�_F�𴆶�k��k3�O�����߅��>�ҁ�W���R�	�.��Y�g[�����UȘ�.�����hc��P�l��X�e����c��C�s_�/�E�a��+���+�!�;�C1r���k��)���A�Ns婸���$��>i��]0�>�k�ۤ�P���:��n�Q}�vb�7���6��n�p���G�GU��r��	��~/�<�!�H��'rB��D�C2K(M�۬����g�E��(c����T�z���� ���Yt���
����l���T�i�$�A|��z���p{s��	������#�˯5�LPT:���6��t���a�~�B�yN�=P$��|��������=S��O���,����H������Tw�|�͆��^��$f���$X�虪��[��
�'9k�]3�5��y�r̺v�o8�:��an fy���ZB�[������o��@����&���>7����1��7�uX"�2+0��wi^������kX��!��5�.�A��������p�s<��ЮO�^�(�a�:����^� �^>m�s���>��w��^V�ȗV�����^�D�� ��U�m��G��1�K��s��o��׿�����&��xQBpG�����*D!㧍����C�߳]�����U�՟7���������	��1�|g���|��A,�UU5`���ul<?�V�>�N��_A����̤�M����Ϧ��?)s�s�>�)Z�gq�=�=8d��)��?sL��H���e��yc������0�E�k ���(�ʢN�0��N�����_4�1�.�6A�H�K��Ԟ5�i>�Z�o�`�~[�� ���d�[}l/m�[}�>�����v������"�@�ît;F��y� fO1"���q��Q�/�a̹rʏ�e(�b��x��Z�[���$�@�B�$�f�ڠ�>�N1e�#�����w��mH}��*���B��/-��R%[4��.�ϧ6���GIݭ���n�.{����?��-�����i���)~P���T~_K��g"@�9}��߅޽2��ƽؘ=i`��o�1m�;�[�Ы|;��Y��^s�=[�9�z}�:���6P/S��u�w?�۾�O�\N��w�O�շ����}��o?�9�Ν�o�ocsw�?)���5�so�!�c_�@ɯe��؁��>�BSg�!�ƀo@w�o[����d��ͽ���]�=�8a�0%)��������ܨ8h�ζ/�B?��%)Λ����o�٩h�k���KxL<1���&���g/�i4�lFw�_e�^�¾'��סOI/KCﵽ��Z����R��r� =��N��'?é1�)'�L|�b�ܮ77�aM���]l�ڣ�\.������|�H�)A���ui� ��i�����FY���Ւ�{�T^�Ϗ+�e ���r�U������s9�����i�᥌��2Ve��ҧ��
O}7�7Ϗ����������eMF�eM�ȊE������hqHM��2�4�*�x����y�`��(��&i�򿎟jêfP�lDqea{�X���/&��)>$y���p��0��9�W��4y�W���*�?�@�j�Ȃy�ـ��t@��m��C�����'`�����[ȇ�yN�U���z岪�C`w��}�N7 �	Rߧ�+y�"�;��5��Xd��4��mmK��հ����D@c��:�/�<�HWV���e�M�����t�k�Z���e�����Q�=R\����h�Z�:zq[˻N�[�������1���ɋ�p~фkݩΞf��j;�������gq�_��a���`_dO
ʤז?��	zf���m���턬����=���H�)��_��}�)Z��r�����oW��p����q�|]�M���SV��ŕ��(0dlZf��ёPq�//EV�BǤ��O����U��j����:�0K-U鍿�G�n��qL�sGӢ�x҂�g�|�o�[9;0��V?ه�&^�5rS}�l�{P|:D*�4��K����t�rR��e{xu�p��Ѹ��UB{���A�_錍2�^���+=h�s�jn@J���r�Zl��4/�]}���%�p޸���nnqW�4��1�Q?��en�N*L$�1�ɫu�H��e���0��`����pf�v;��6�{:�G2��hPc�,���P}q�6ßBZMZ�$��
n>o4��k��ꭥ:�#\�:�����z###��%;�#�B�5����oa�/�����;�g�nd�U�7 Jɹ����c܈�q��o>��6��[�Ͻ,���g���a��/�ţ���W3^��}���'�7��2��=�s�L���[�:�0]1k�6��J񺼰}[�{��e�N�1���U�9L�fCv�����}0�W�\����"�<�~K��b�`Z�:G�4l�F�XK(���>�+	L����d·�- ��oΛ�7@�6�|������w�U���*h�E�ĕR�z��������e��
������k���N�l5���)�/�m%a��V�H��sE�k�L�L-�'K�!���MA��'�s�?�`��A�8� N��)��
�'�G���9��G����|<�'�ـy�|.P� h�c8(~���y�� %�y��l��|�<g�u�g���u`xԏ�6�"z�3(t���!�2�͙:�� ����$�B^!Q���z�4�O\md�B�!�{�d�������" �$j�ڿ�&���u}(�nK��J��$��	�	�	>D:Ċ��ax�rQ&,�,�,��@�h�n/.�&�}����~�Fڛ��VV�¥���B�!��@7`�`����ܤR��� �M��������Ɲ�qƷE��D2Qҳ�3����7�:0����ƁǍƕ�R�(ɦ$�p�`�Ehӷ���2X0��Z�Y�m}[���)�fV�2]�KSmG�vы�tt4�(�lZ�����k5Wϵy�D}��W7�����i]�������5�V,Z�W7�3{\����ǉ�$&3�22{�ɬ8�-*�x�Fw���jM9�f���29E8�nmC�����c�xdeQx�R]���Q�e��>�xQҭ>3�-�2ȣ����2�a�����~������O�²��쩍��q�h�)1=q�X������������������=E��\��߶����h���=H/�L�g��;	�i�WOd�+$r4�ߵxG��D񍈭n�J�ò����mBSQ���X�� ����`����@��@��8!��S������.����b�g�.t%��7������b���mW�����R�S�Xm%����s�{0{d{{�{=�K�� e �e���s `�K�I����	t	<M� � � u���Ă�����!�rt�v<��.�v`�UyiErf\7�y>��ͥ�0�ɔ}C&��6@٪�hjN.�(`�m���T�Rמ�����g�w�^诠xE�eJKLe_�L�I3-lH�C�h΄]G��f_{�I=]����z����L�[��kً�;a��IQ0�^E�?u�7r���>h���w��mt���.Kt�{u� ��q;����z��S��GLCт�CN�� n���%@���&��dd�x�F�Y!UDwB%^a3�l^�|�v����4܀W�d�W������j��[Y\����	8��7٦�'���K��=�����|�g5\i4�c��/�}��Y��7_�tw��&��8J�HjW�A�k��W�UZzK�+є��|*��W��'Mg���������J�9����_�a6��Y��e=K��C�7�̪�ѳ����3X�����5�Z�]�B�0þH��;|X4��u��)��"X�R�������#]5�w�_\����y �u�R����zS��&��O��Uهçz�s�ݞ�����K`�o�ȱ�9�!y�����$��b�w�K�eo;�J��!��B'V2��A�/t�:A�s���k���瓹�-�w!S#%�+�d�0ʤ]�K��׍�Hrs6�9��޹�;~ʋ����.��ň��}��7]�A~��=�w��]�(�7��[d�9�f�\,��O��4�ވ剈;a��P)q��o������7͂�l��:��/V �t���ǭH�#�a+�'j�*����A�⫡��U[�s�u��pv��Wo�P7���Cq��i4xi��,���`S4�z�(������Gm�ۊϚأ�/K�(�]�5�Gy	ϟ��s����=��׾DV߁bŜޙS4/���ħ��g�WF��Q]���zof��~�߁����I�CJ�*	�,������ɷ���������mi>�����8�,RY���3�<O��&�0r	1��H 4�����.}}��y��y�7��{)�mR7�#�=z�V�R���9��P����紿o1JK�2�r���Wd�,(Ь�ܬ���-�j0'Q����Y#K�-�~E>���=\�y����R_�����$d[��t"1Pf��w1	,6)�=%��	2�o�|�Z��J9���H�UŲs��U��J�9�Mv�~{)�m���x�%�|�Y'���9I����y�8�������<p���^���j��6����}��ݖ̱�2���͗����>�~Y���>5�����*>K<��9/�{4���*fc,�����
��m����4,U��W�*no�?!��Wh�C�~����n^*R�8F�v8w�R�w�zfٿ���ni|͟����]��C2o �e�[���z��m�MN�#�;���v���2��'��P�#|��Kmd�.���%��~��O�tl�0��6)���K�J�u�2��N򜡙���;�4V���V(?���~��}�x�祫���L�i��1�k)Y&Ϲmo�Å��LaK���N��^�f-�m|E$��ZT(SH���.���##ǆ�z��3ZS�b����[�M�h��3GP���������6�'��ǔ��,���!?ai#��("��x���8c��Mj��
F1͍8���
;�X�x*�9�Uk̒9�[�3�.�4-@P>��v(��	lh#�F��&�S�$�N����l��aJuM��@쓡�_(�L�3^�'�6Ck\�wI�]SwH9����_�L(�G���h�\OA�T�_�3�a�� �~C�zX.]�P��1�|H&$,Ε�����.,X����z�"���S�]^կ���$6=:e�~t��0����v�:�I�����t���~|�q�þ5��?0�����oq�1W�#���v�Ci&�Y�w~#�������}�fY�U�=V���FX����uޜ�{��_��ֶ_�=�7���j��O�G|;�<�&��F���sZTc�.�m�s��Z��Kb->��|G�ψ|��$����'Q� �d�FYg�z�y��#5C~G̈l�	� d�`B�r0�ƖK����/�_ܕ�3ϗ߹�_!N",�i�T�� �~�=G�;Q�0 ������0D��\�jT~D��<H<�JĻ���
/*��B/�����s��m�9�g��G�i�������>��W�4u�iߟD9���k��
��T��3f�y^v���`���y&>'t�ɿ̲��0�Ƕ�ж7@qkrQ���#���<̰�6���̖	�v/�5
��N/Xl����T{)z6�v�Y�I��S�	��u�σG���"߶uv�~�Zv��	�+�Y>��S��2E|c��Ɯܻ)Z\L��/fx;3�;�����M�$�.'eL��-'��_s�UP6e�'�'u������ݓ���J��a�!u)�&E���F�����Yy�~�g?�Uh�VK�x]*�z%�{�
r�c��D� �	�|�\���Z�ReJ�H�o�)��t�/�0�!}����=3��ܵ/���q|�Y�D��� 2�9�"�ڪjf `�z�:9o[\4�J��}6ٟY�Xv�o�)�i��*�ƴq����-w��.$��N���V�->Ne��ޕG�j����!��p���%�H2�F�pr:�M3��ϖW�T+�&���ɰu��y�EY~L
�nAgqɴX���kY�>���K���- 	D�v�ro�]����5˫�h6�*��Vj�,;�z��!�w�ŏ�~���,|�;u�J��ۻ?������޿�*[d��į�oZ$@��t(��}�r��hF���ӬH%�Nq�4�yc �0��:�Ͼ!��x��%j�WW�َr.	��]��|*�Q��G�Y}&0����O#Yb�T�_�0K�@��t�r���q���_��z]�ׂ�~ �����d���������{S;��ৣ_:_�^v�����*XWh+|�ۭ֍cI {���`�����b3��3�e&�̵}\�_�(��w�u�q3��
 ����g��
xie�0�:۰ ��F��g���/�ᇗ��n��'S�)o�aX����q�)�ͺ@�KC="k7�g�	��pY�8�x�Y����x� 1-��O�H��x����Rej^�q���F8�N�����_�H3"���Zӵ(v<#}�!��[�ԧ��a��Fx�N�_zX��0!D_A2�u�#|�W�V}�-7���2��Ny��ט��Ũk\ M �/�9�1Ƿ���)��<Cn#�1��jN��2㣘�q�lh�-��Bt#|	��.����Z�^v��4�@��~�q=�!ȫ��-Dt�B_Wn6#sz%���)�}3���ߌ���-8֌h���>�|-
;��>y�G׈H���R �m���(�A{��R�;�,��y�Vk{K��w���35���߀(��Y�jJ��20ዓ��ɕ7z�Y����wʕ'Qur��� ���*����?S!�����6��pq�5~R�4v�4�a�2m��2�ޢ�[����B�|��.?m �k#��ޚ�ˠ��1Z����#�f
�r�@�Ǣ����|�d6�r��_��^�=���ʴ��s>q/�@�j0���M��Tp���S��t]�p��1�6h�m@�ML�0�fl-/��|rsr��a���Tt�Xc���Fj]��d��-�����i�Ӿ�!x�+ ��\R�)5L�*t�i�t������:�c���%���nI;�����4v⮾�)��x�E���۾?.yhLI(��]t\��CC(/�icC�.�Pж)���.��d�V��n��HX�W-��b:�����?��{�������[UU��K�|Gk�.�Z�{����"S�ea�ydO� �p�w
��/�ؿ�UT���K��QD��Æu��������q^���6�sǷ/�cǗ�Ƃv/�_�ݱIl���w���}ͧ��ئ�癛!���H�P��� p�;�A�[�3gl͉Y�3k��-����,P�7Hq6�7�x����;������9�}�����b��sr?�������(v�;*9���;��@��y�^�,]j��]$]��U��BL�7�L�3�?������w�����P����B����a^Uz���6j��D�S�I��~��,Q����BT�����&�%�қN179��.�D�j�m7E
7Lۘ[�y�~�~��-���~d�3Qi*`{`�6��=�y؋t��c��͟K�		~F���Ɣ#4C:&TM[����*!�'=�|P$�bԀ�~ܭ��4GW�F♴�n��F���hf�H<c� ���,_��ϴ/4����'�#��ɋ$�ڍ�?G���,Z�K���ڤՀ��w�g�%�,�akֶO�何��Ϙ��G;�-Ƹ�\�V�����{��ȯ�[����n�vX���#�~����@�#�\�dЁ��ppw�ꭊ.�T�빺�>�k �`��.�'b�9�T@l���#�eT��+�`��!��	��)��K(ٿ�����g�V�_�$�c�E��K;� H"��/�7��7�!�A�l"c�ْ���. �J�Á��׎mb�>�O�,C}���,ɇn0E��b���#0�L�zڇ�('�����ɨ�� Zb��a诶�l���mډ!j%P�뤣�~���<�/V�(�c_�i��c��h�S��O�窞��VF=;�΍^�6����k����?גv
�Q�]�l�=f{�����g�p;�Ǽ�Z�j~�=D�{���?�+�i�����;�Q�n|���r�T�o</&�N���Cݻ�r�X�ݻ���Aci��gJs5�	��/�IO��
���"@̈́J`&���'1;U:�1� �K�J��\��	 Ѐ�~1C��n�d��ϟ 4ѸYG�:S��j_xd��l<\�*�m�(ؤxX��Q�}�E��\_Tx���aOQO����0M=�ZN��?A�t��F�ȭ�T�� v磃�8Rɝ�����1�t����_q����x�k�=e�8���0��nBb��!I{�R�ݓA���-��]վ���%���\�[i����W��
�Ĳ]T�ұ"��XS���O��sM4�>E��Η��W�Ċ�<��\I���\B�\���9�뾄�
!�=/�D�@�E��'���T��wT�{�=�=�;zG|O �C�����]²������)�o����_:�>��a���o��Rx��������@�����[�G�������� ����_D��O��.�#ei��3�3�|(���ޟaFK�s�Z�W��%�|�y�3�a рi�Y�_jF�
2;��{���ʏQ��J+UX��+��D���c�I��ۡh/�PӏrDƓ!~��%]p��3(#�	���L�	WU]�ؓM��%�.����n���'ϋ�TǤ(��2/m��U�;�;�~d_���@�����~���g�@z=������^�����n2�t�?�g��Tk���-��������t���ʓ�j�И��$x�
t�zq�9�����պ�)>ĉ�\S����k��ER����<�ߓez+Q`��Ō��`�'&��-����,����n�������+|�}�r5}f|�o��O{�IO��Z\,Y�'P>��(����ԁ�(2�݂���W�vY�`y�9~}��Lp ��Q��e�n�����ɳ���j����B >�,�>wSxC�G�B�v�-��甥�E<=��]v7�-�=��
_xM��{��$�i�X�N;|���V4WLw9M���?l>5 Dt>������xa��^���v��/�ш�S���Ch�w���sӍ�t?x�G>N�{��h��i������4f�Ml�o�>z�� D���szkXz��w�ݖ�~|����W����?we��p�w4���Zn�k�I�v�,�Y��+BLC�p�+�Me�͊�I3`��|�¥�.��\���Ɏ��4�$�|	�!�F/�nCO723����>�zazq��g����`�u��g�<U�i�j�_�i�z8`�=�B5{�p��f���#B�� B԰�3P� ��&��}&���� �	��|�e�nS�3�\,u�A=}	�������z���Vc���!`���K�d�]`�����y��o�B�w�H~�M}��}Z�y&_ਇk����gB{����f_���O,��z͍����6�	���'�/�N/����Z���{\�]�<oS���ÆF��W׻��q�{�Ԗz3�'�S ����/2M)ߤ����%V�|:[�n�OQ:A�m�� ���7�}ޟ걽���iK��w�1�36}��#����D�ުJ..����JU83L(V���p���X�/Q�y��pIli˾�B��}���iVy�~��K��\���~����H0e(>��a!�Z�����	��|l����ܠE�:��*aN:��E�x�L�v�o��h�.ސ�Td�5_�"�gy�Fy�1g,��H��/��_�%D�6�H���c�}����t题��ķ�IO��#�E�C���Y�X�Y�g�e��?�u�	4�l�čd���(�@V�N�����t�����=?:��@�8ɸ�=_�\N-����Y3�>R��{�H��t�?�&�x*<�<t�U1�W(��P]9��X��j |��ix���H-Ya�TK�J��^���\�ɋ��9#�S���E%��ǖ|g��_�쩧�<����̼ϡ�}��rM��ʠǻ�������dK��ee/�� ����c���
�����aO�H�R�O���F4�}�)$uQ�XbG2���o���o�|,������c?N(��i��{��G��{�a��d���a�3�(w��M��k�k�8\\Y����R��t�����"8���ܝl /��?h=�^(!�Ag�}�S�f��ŻJ��૤�bR�N���)��������ᬯ��U�><s�*�m�ޟ%����r���d�c�}�"�UXDY[Ӟ;Ye���%�nDBJ��ZL}\qv�dAz�S�?G�'�S�*�mK���~���߃�O�͒�i���>���i��W� ��\Lnz��u�-���ۇ�[J/e�AP�\���l�m~��`i��h��6'��/��[���t�XIU��=�� AM ������Z^!����?mU�6n
�&Wl�3y5�1ߝ���햕�-�rz�9�SEQ6�W���#nW�Ԋf���O)i��_�M��E^��"�kt��?c���ԭ�MT(�$�b}vS�����^��d��W�W ��	�@B�]�V�!��_�\��A�Q�`�/�QA�;p�EC�_�~��=X��k�9P<�v{��uh$���]Փ)Q	:�6��q���S~<6>³�����Ԥ�l�kr`P��+�T��aWŸ�tўs��"�U��|���0a?�S`a4� ��K`g�j���>�7��$ E�n�zh����߲����G�ߺ�oO)7�]E�
oȺ�rƉ���sj�$�������<��&w���x��b�`�����K*uT��\�n���v'_���R�zE������+\�'c���(K�F�NۊPe�K�*��T��3��'�̻�dG�C��F�ݰ�>>��{��͈��{��3����C������1~�� �娃4�5�P��EĞ~H���?���l�[n����D%&��6y�'�&�"D!� D,.����|�o���4������=�H����7N~�:����m��a��y(�������}�����c�D��}��2)����E��������]Y�LI��l���������YY�\Z��б���>`���Ɨ-p�~�aY���Pa{�!K����%?��N<��&�����ۀLs��GSx�K�τ��~,%�x��&-MQ��*�Z;�����ogⱘWļƯ�[����ч�A�9אi�6���<����D�����H�5&�^�vs0+�=i��88�p��Mq�5$���0W�����&���z���#}�5����JV���$��t��3�9��Jm4�����w-s�!��߳h +��*�ɼ��ك��?"��|��#��|er�<Ǳ��ff��H�rX:_d�'�OP�Y����I$�x���Np�v�U��u9�S��`a*��_�L���T~?	mă�2�	1Z�6����(����+��='d�����(6�t�fR����p�3Q�O8x���Y�~�)�[�~���ɺlԁb�65��x��|�q��MH��J�6!��#����;��˄X�=-y�Y��) ��z����MZz�t�)�OJʖ:%�]=Jv���RHb�@��'֟d�9�'�	q):�T̺�i�{�؜J懚��TR!õ���c$_�
8+hN�N�ٷ��g��O������W���u��S|�c�%��'(�<��Uܖ��(��֓�FP̿��yr�ab�'�)�������gU���s#|�.�J|9�v���\O�_�<��<������+���py|h��z�)�h��@{�Jҟ�L|��d�-y�����^9��X�r�@���w��N���&�-�+��-²�E�nɱ:��EA_���kM��;f�>���}X�w'�}ˠR V@g+��/��>yr2Ӕ��oǋ��+7�7A@#�p��`
��S}^��;��!���P��O��%����f��)�W�G6v��qϯ1.�R�wNt�5��s&.o�>դ`R���]~Q����>`��OQ�1?E�TBnt
���U��&�������9;޺G�l3���SL|C�Y��+�3Q�V��E����X�:�?��:�C,�7l??��:��|�e�{{��nE؎�4�߶�����﵌Ԛ�~�E}Y�Ӏ��-T��w&+����]�>��o}&����c*B�1w������.7D�Q��#'�f��R۽�eQ޸��:[H]�HJ3K�{z3 ����b,b���`~����N�.���Y����}��!>�����1H�p'ڸh�ո��ы��Ζj�]ۻ�1p�;������~s�H�����8X������I�{܆z琈K�kB\�'۵���,\0̥���ckD]/Y�XB�U�|�A��Y�hy�gx|��UfsI�}�yi��9z��cױo<��M��CX�sm�����d�{�#����f3���)��h�����*�����<�v��h'��ܛ��cy�9�Ϻ~����稍��=1�N���>��~�?��.'� �����X��~?x�Jv�BF?�0P�_�iA��u�������
��tO`��N�C;퐉�bD�����jNGtsҧZ�Zn��I	V[X��e�}n��jkЀnG��_#���t+�5h�_��w%���%��t̅�}@�F^V��<!����41C�S����>0PD�E�$p�wĨ���I�1�l����¥���TCX��H0C��"�PmI����x2.��a~l	:�!�O����0@vd���QD���nx/���_��D?Q"�@��x8�z@h5�>�W>Ζ��ޕ���\���R�d*�匁�T����BM��S<Q)������܉� Ku��Hȃq���F�{�T��ǂ9�$ϐݐyb\A|�c����S��!gK:����Qx���˺�1��.����H@Q��S�������Y�AU���F�\�2�@^�uڔ '~�y��[ř�9�JR7ƙ�j!�TaHn���?B���q�E^��H;�0R<��,
9�p�z�TSx�ԑ?i@���B��8��GF�n�'���@	H;NtE��A�cm�!��0$��ł��fK;b�Bc@��9�̀�!�g"��sӞ.T����{�`�$oAyDo`}�o5$����H�
�){�AYP��w�J��
�Y�I8�ġ>�_���������X)���g'�+7J�h�<	�B��#ِx4��Y�8Y�ќ &s=������gZ��Ə�����`7\k�P���B+����\&[p�<[q�;�h1�V&B�5� ��Z�/E��Hޟ^'��Qc>+�$}�L.�vz��D:e�M�T��MQwo�k��%�"��\&�k/3<�	��ʤ�/�d8ю��8� ���$�1�^+|����
���r�%�4�&�(������qN$��չpټ4b����Vi��6y���z�dxÿ��u˘�^�@7�bX��뗈�0��5Xo�_D���>��)Q��v�rKb1q/n�U�m������G��G���)��DJ��-��݄��De#n�f�=N�֒U��5ߔ 穅 ��s�/'��f��S��t�徘�	�֠��$J�3�}#�j�����8�G	��\ɛ��G��/b{d�`��B�y>U�`�<)��,��%��@���"87��bp�e����i�n���7:A��J4ƞk�̣���B���L�Ԍ���i��]�� S�la�[6�̞���z��PQ|��h%Ñ��������5�K3qZJm��J��k���Bv����U��Lr�Bv�f��,7�Ugn�=��3�I�&7fu����Nހb��w�-�?o�GʹnC�
�T��'r��PR<vʾ--T׻�gQ#n�����D���_A"��ټ�:MX>g��u=��
ټ��+�iO7�:���Ů�����[eQ[͈1�Aݛ^Wꒊ�Ed8&qZ����T�q0������R�ێ�8_�	5��&�s��\v�!���Н���mj�*��ZL�	��	�&!���,:�A��
0��P=��h�!2��By(Х�k"ɮ6��U��3XXV{�2�|f6v���b�H�ʹ��@mjl;`�5&9���W'�9i�ܵ9�2""1�����і�J%�7�l�z�
J�bD��&�Y-�xf�ַ�`��l����,;0��Oދ�wb(��3Оd�H�`ny̓iD@���o�;�H��r<Apch�}�)�k%.h�K�~���:�>���r��aY������Wp���<K3qi�K��(�W�K���fB�u��{[�M�����d{V�Nm�j�tޗ�t�ʎ���̝߻,s"h��S�v�M���J�^�)I�O�A�)~(TVh�S��/%��~a���'��)���6>�l�T"_�|��bU[���\�>Kq���	�AԀ���N�M���(�92�'G� m�3� }:�?a�p��˦hi���M�D���K��Ժ���ƲI%l� _<x�,���̛�=��8�5(�6p��KJeˍ"�3t:�W�ga���[��4�<"���*+�k�'���������O�p���l9M�&kW��9��4ί+ܶ�	��A���w��mU�[,���B2'*YD�O]j�|E�嵁��37���ii6�W@f0�Nq�Z{��T�����ܢ���Wz��qώ���j�Hy1i�je�iq ��܍�HL�HS�j�a�i����y�v&7��ZI[��vDO�e 
���`�w�ͽ���@��˖�V\dx�T�V�Ya%Qf~�W*�W��&�R\CU����Y����G��P}B�9���ö3w����Y�&L�����%�.���Q�I��B���
����E��+Gu8̯����8�	����7g�lp!Jw��i��1,pުnP2�)(�l�}��G�����ʶ|���EZ�.\�f���x��b���r����c'�ӥ�x����k���@�T#�ڕ�Rŧфp��\;�TLi���jRQ]m���g����Qo�����HF����>��F#n�=��O�ó��z�,����2�~^�˲�pd�
4ԝNCT�6ޕ*o%C�2�//U=����D3�"����u֯Q��.9�\�����t5iG����8*ԻT������p5����!RRx|z ��v�M-�j���	���8,��	�g����[���/9*t��ô��ɍ� y� �Op���a��}zPx�8��O�;�W��-4Z��7�f��h������A��^�cҝC�.>��t6����1�5��N�Qa����AT�%�п���� )u����j���ݬ��^ط9��#"L ��K"E����I��Pg9�f2�6n���	��gWKDOM��h3	��8�_LP� ����?�9a�\�Dn�@i�V��fx������E,�e��]�{樐ה�	���>��\W�7�wݥD�������?�u�8�?�<�,�\EjD*�=W��O�/ai�����0�����_}�~�9*ys/��m9�0>ղ�4�*5)9b���A�( V"�**X�S�D
�kUe�ZL�a9Gي�)�P����
C�p��C�D���3�2�p�?�ws��n�xI��T�{=v?w^��v_߻}ns����`��J���Y�������F�[H	�n��59΂�l��T��ˎ񞺜\�M��&��ɢ(��S�$�x�=Q�مg����|>|J��%��_�2�y�~=�O�ET������'�fB-�|�i"}������]�@�٩t�[��
h��&�p�� ��K����'4K�e���A���gY���$�sH����l�ܰ�-H0?-�_�Qѫ��MC�x:�Y�I����?\'y�\�4D&E�� %�p����%b�P�(�V�>��o�!���@�r|;�1���Ѵ'��.B��,`�m����T�0�Fe��B�\iü��/W�go�R��TŤ��B%h���a���w<�>�Y���<�:�Yd����-���~����F�M��-u|3�3���%�8��ϰ��.:�<��7��Z;M���_�~P�1h�2�,�3��B�_?'��n�n�k=��{MK��n�{�����5բq�>ǙJm���Q��o�l��I1��PB�:6�Ư�e�]-�εϛ�ׯ=�+Av1�n�����������|��k�:�#�9���*�.?�Qp���Ʌ���{�d���ۓcL>r�k�p�*�A~�����P���҇���*�B���r���k�J�|_!�B���A�j_ލ}Z�)wLW�,Π,?ń�ț��#-�x���/����Ea4�Ov^`a	z���w��*�?�	j�c�9�
��&���&�����1���o�哠lkj|�~�	���p��u5r)�<�V�R�*��;��h}�s���1�H�'�U��G�ւ��؛�+B��K�����9 �p�v<�}���o�V�|�i�i]پoїqؽ��q�'��B��p�V\L��'�n��eV��������ш�S?�@��j�}���@�@.�J�F�D)�U� �D�NhQ
7t�?v<M�{�u¯삢~1�N��;s�g��{=�k���3��Uř�0:S�h(~�.y��)�W�|��H,S�m{Yj��*N��(b�T���_w���\C��7��v�d}[���h�׳ud��l�М?��O�%�D�D �����o�Ȣ52�GBgd��Z��,�����
�5�
��.�c�A
�[<�"�Iz��S�q~ߕO�!��1r(���=�2�Ȳ��U��s3~<ֽQ��'(~>�#�_����1�'�}x��=�E�-�iz�+�p��w�����O��R��I��e���d	�bL�ۮGl$����:��ٛ����%���1](%5��W�*�.b0��y4Jp?���k�@nQ� b��P +�U>�*(��[.�4-�O;�'��`'H������+��p�����I{:������+�9�����;�����G�&���l	�,�X
և������_^���+Z�0\9��-�( ��;���>��4Z\��Sr�2��Wb�zx
��(����t�v�Vǡ�w���9S��*P�(:�*Ʃ����W�k�d�l���+��������W��ЭM& ����v�ٟ_I ���1�R��1�q�ɟȜ'��y����L�e�0x��I�bT�ʷ�M��_:�ձ��05��$Q�����߼�n�
,�72<����x���;-�3_q��T�!�C���s�m�5�Q��+��h;`u]�yh�B��7�0�b�����pS'y'�Oߟ�t{���{��|�N���n���'��O�C8pD�3�~ 
x���YP˕=R�ąt���<��r�Ս�vؗ�Zx�a�̤�_J�<��*n<2���b]f;����'[�3�h�0QY,��g�0c�.;mh�͋��~s����* 'x���E���t�D�o}e��+�w�3,��t.͈n_Q^���O�"�b�
� �. �E_|s�����#��t��J^y�p�Q��A�B��Ȝ��ݥ�k���p_�b����Ocqх3T�s�{���@syYa��j�'a8��D��C�Aָ��jg|��OZ/~(kW��`�vW$���
*�?���U��$��F�+=^�>ʙ�����z�M#�O<D>̳�,|��:D~�d<�D3��a<mC��:�]Ґ��駋�%��n��7�'D��Di#z�KJjX}�� J@ �DO奜.h0��0�=�vu��}'R�I�8�a����Ӈx��Ɨ���z)�5����6�Pĺp��0��n�{�{�jZV��(y�Z�k^>=n��.`ϝh����W۝� #����?($F��S"il�Ѕ�c��P��$��dH��u_�P��F7��D/!Ƒ���QC�1��z��8&�8V�ҧy�ύ���[�T(��^Bo2ȵfpY�I��[ܘ��F���/��8��7MP�\�U5*�N�msnY;�J��AA��&U�x5�$��d�X�L�ì��@�K� �PD�4������l�ᅽ��a.V]���ަd o�J߆;WD��n����d^�n�!��A��"̰��B�9�.8���1�u�*ˢEQE����U�=�J?A7����5����<C�1��u�Z�����������@@���������%��bS�se��V׈���nˠ����,ͷ5���'Tk�Xt~��5F��ا���$E1���b�r��aa��Ɇ��ɇ$��g�6]�jw�(j�/{��U�Y���$��%n;OU�G��Ӭ�Y��r���;5��u��`�uxF�q�w�.�����\6\o�Ţ��o��N���@҇L�g^�gK �0�j2I	A�}���X�c���G��_���ӻ��H-{�BU�֘a$$�b%T�:�1��:b�Z�[|ܗ�O
]��f���Ed� Ie��Y@�W��;&5���P���@�q���H����q�a��w�[^�-���V���D8�X���:�`�h��Yg�wO��wz�?�4e�#�}X���H�>etw�����*G�/�U;I�t�Q�&-�LɆ���D�p�v���!0;���?X7ѷ��q�{�Y���[�}kˆ�M�QӴ���K�`�z���7t�=<�����yEc'���"���e�*���t��f�j.-Nw�?��s�޲_�������o�Wi��c�K��7�����i�����U]0�1���nq�W�7��ߖ�?�w�/�S�*1lg�:,}�׸����_o�F��KȔ�xOV�P��a�rA����M�)\�b�ܑ�G�Kt�]�y�ܲ��j�x�T��ϛ��<�V:�n�)��A
�ɰ�D��!����H"@d�j3`¨X�C0.�����c��@��G��j����&�MD7�DJ�3
�r�e%��p�����x��}��m�}�����~�z���;ը)�ח���@�m�L���w��q`�Ɂ|6&�S�ˢ�I�b����"W���
�5��ӳWP*�\��V�dA}:�U���Q��[�E/[���8�Q^���|���6��
�!Һntq++��c�3~�l� _.��'%u�(8�[���AD1/%��#ќ�H��p}�=1ۇ�'�xb��7e��.������Ch��i��H�^�&���W�3{��B�Aha�ث�6V� +Z���B~���*�F�R�A��=d�i����������MM�#��]Q�%�𱅆Hd�L�.��1���T�&$=3���#�Idß��d=}R� ���7�'J����+���h�[�_��G�����`<�/�����l<�ϴ�>W�����k���&�;lǛ9ϋ:~��QT�5��ȳFD\��A�З�2`{�~M���#�/��������������v������4��j�I�^�?[�}���l��Kg:D�p��q!��Ӵ��#/�Iά9�RaA�dU�S�JN��o��9t��CW�l$>��f$ ��EL�Vj�2�k��H/�քÊ}Bſ��Ǽ3�:�GE�iY�ŘS�N'��G�㰟�1��?u�����d�>w�-o��>��i3x�f�ռ����8ܺk���&��uO���(k!H���R��G=����c������Teq�°�&9M��0���S$1�\�����bvȕ��m�?��5�a3��lnk>Z�8v|�*|��"�� !h����Qܟ�xG��OV��[�Q	$�J��3��Uy���Q�
5��'F �9 �@o܆{�k@f�'���+_Ti%��w4n�<��nݝ����g�5�#���?�\7��Z��S�x=au�?�tq���z|~$qY�y��ci��K�K{����Qe���e�e���@x��h���B�S���uj���������������&��;�x�i�)%������i;��E����W��i�!F` 4�I \ P��]����y�#F��$�:>B�J���m�-i�FHZ��N�O�te�U�U�k�ԑ�[��=�*}ZE�L��G�!���1�y��n)�-���-DZ�k���˺�\�L���KN�k-�n�Uu�A���yۇ@��7Ӟg��7�o.��wN� ������滋_Fm��B�7�D�Ij��M�Z��0�G�K����
-�z�wI��1���w�(v�G^k���� �7��!s>V���.�:�:y��D^�onί�՜�%��Jp�b�C���w� ����9B��d��c���$�A�p�X�B c����/���=����(r��F��@��f��M�b��/?�/���$���8�?��7Ǉ{��=�gd	�NS�e��<������z��&}�m��0;��2��w��Fg�B�p��T+���r�M�(�Y�e^^!~-�kb��Ib#[�������5�<�Ni��m�l�Im�#ZDٷ,W�j�g���݆\��~<8�wu���d�Z凪��u_�?�f^.r_.���sz�Y#Y�X0ѹ#���8���x�n�Sa�i��K8�g0��� ?l�� ُ�����},r������:�z��aE��zW�`�8�l榅2���X&�i�}0iq�h����x�7~�'o��7����c]��r���!:�����_v;���?v��������H�c.�&�����H:�cؕ��2����=�O+/���E�
�|K�+NQ[�r.5����)]2c�d���\�����$�&����N�Am�AYtG���_z�'�[�W}M/~=��ݟ�Ŕa�a�^F<3Sc\�{g�=zg�)�Ǳj6� �LT�b.=�?6�W���B���=Q�.�=�xN?�x-��E��a P�/���wS׌�Q�%ݱ Q��F_�~��(}<�t��)��\
b2��,	з��{VI,�{�Roڻ/��9[��:��T晑��h�`�:6b�-i;�Ї�O�����=:�bm���$��v�vm����������I ��o`��*�!X�2g�B[��y�ת�k����w�ȝ��fЁ�����i�W0慶-x��?c}0�W��
O��:��Gw��,��?y�ʹ!��Y7��.������'I�0��s�Y ��g˭�W'�.�R�����ږ�gɶ������7r�Awwxg��7�8>���3|��o��(�T.��u�=Z����C\�j#?���EۛM�G��p��^���Ar�mr[�����%w��
|j��j�_��}��2� A��?�R ���`;�V�K_�}�r�+r�ursM��>�iV�g��Ѻ�^�y�In;�`7�:���Q�f�P���a�%Gq�ˏ%�@�|^lv�����~K�f&��?h��ҙ�8�q��O��8���Ù<8���>���s�z�W�tW{b��$��_�"43҆M�v�0���KQg��W!�~$!C:CCC`C��;�oOӁ/_����]��S��O�ˇG��_y���ޜ�۵������e��Ǿ����鹾�C3��ί/��QoS�^�����<���-�����-��m~wƋ��Mɫc�����t,� E�:+��i���~�x�tU����+"=ޯ�R��鹓'�lp�'	���?\�~lC���������d3���/�V���m%f�o�
 И�F�D�C0���q�����OZ`���rF�6��-NDGhx�n���o�����K�{]���(��^�[a*�'�TJ��ʓfE�U�Ѫ~Z�z����hK���;m��'R�f�C������a�l��z�I������&�J�\��;{���lU�%V���eD�T9�ĺ&b�N�\���9���QҸң��0�{�>�+�f`ǎ5 k�oA׎S� ���oD�ouTT[dY�������|gZ��	6P��
�B��Ԍ���c�gh�� o!X� �K�v|& GAC6C>C��Go���3A.=vP��_{��>�'�l�Oi�]j^��l��X�]��[�����+4��q`�;�t�m�ի8G�l�w{�U���vS!r�=��k�׻�7n��w�|[�K��W��������o�~ġ�W�v/ܘ�;��m�����|W@G�_�pO�0z�z��_�0&�(oC�Bo��-�]���
 %��d��j�2��s�@T�5@J�ld\V�̝z-ŏ�l��D��I����a{�im�3L$�j��Hk��F	J���� J��ߏܯ��0�
\,0{|fR�@xV�����^��t��u:���	�v.­@H��v��ĞVQ�W����SG�Q�湇,##������fޞ�
��`K�5\~�2�،�:�Y�v'�ǰA	��!q�n