kV��<T-m��.V(C�����GyG0��݌Sa �!���K�n�s/�i��b�A��DS(G{
�����⃇��j����� T����'��<QUQÓ<��`;~PW�1�N���c�e	��T�jX�6?,L��7R�� �b�O�Or]��
�L�"���/қ{�����1�?���cf�䵯�K�Q�OX��7R/��hkA���z�~@�V����̠�U�ؤ\����ζ�����k�T���?3���jCsKo�OյeR&�Z�VQ��1�D���I��q��3�d����f����F���Y�Ў����������8���x����;�_�i��A�¢>$�6��5��<I� Y�'��;o̶�����+
>��}�X�>9�3+�&�e'��:4
N!Y\� ��i�z~u��B*8$jL�[�7<��xi�����*�2)�~0KI*DI�5��V��8��>�1P��H�����	::iю�kH�b�r�{��4�P����E]��-n4�	!+��RU��|��#X�����Ǔd��hѱ�C�ܔ���%�Ō�p(�1�:��7	��?q5ަ�"i`ǱI�'�VP�=���u����n��@��I�t�h�=L_HO1���zfl�B���~D8��Z�Doa�
����Z���:��	�e�[x��qLwl���J��3�빊��֖K�߿�}r���=�����J@��	�c)'/�_<�Д�h΀�C��T��1���.�� 0q��߄nثMĺ���`��AE�:}'<'9�BvxE�wX��J�O�O�(�Ct5xK� ��m�h]�a2h��bQ��n�~5&�W�֬/�.�Rm�b驤�d�
��J�9��Y�a�C5�4��RR��|�{_LU\C����vy�^�2-���Fo�qd.8O�����m�!�ױ�+�}����9�ł 9����\���U�aI���/�]��8w%^�(:*�d'
k9���PRW���I�wrGK�Ld�h�@�����"���];�j��5q1]h���i��6��r��h
���*�x,�q1��	�IC]g���)�|�HLq�H�t
�*�s̞��D�ڹ4��~�Zt�.�|�a��C�7�3	�$ֵA(�M$�V_v��k���@ݫ�p�4��?Z[�SV|�o�m�� ��YxD����F��]i��S���Ir�,�����ݶ��3��X}��p�]6����,!_Wٚ��>ɵo@םϐ��� h%��Q�Gh'�<Ea$-T���U_W#�i���Q���%���(��4z�'	S���g~N���E���E�6�
3`�Z�*�WA�ǥ�A�I��M�G�UFn6H���e�YS+�#��������(h@-;1��%�l�i	��T;�\y}�\�3x�\h������q���`����������B�m{~[t?L�F-۳��X��qd��z�q�,MY�r��L���1�9��J��.9M�2	�Z$1:���N{�?
04h��������%-x?A$h�[���#���g6����ٞX7����؄���:�=�FwmڧN���׶n�(�'qy�P��a[P�`O.���a�|p,e�>��=f~{�.J�����þ��Su�'���m4XҠ7� 
v�
̎��}��A�Cud�Վ�� ��6Pq	�]��l�[�z ��4�c���~�Ȯ4��a�q�3e������~�蜽|5�qt��^�M2���������36�l�vk͵�e�Iހ?� ��܆��$�x=���M��(6��^�I7�=�s��ݎ6���U{5�1;zwd��Ѕ�嬽��۵�?�f�Wh�e5k�s�^f��w����eg��`��vՎ^��A���:�a���/#������?ƹ.wؾvk��.�u+�L��6�M	Ʋ���L����sԈ�<r�Y#�F�\���;�:R`%3�c�)��|^�������g�;��/�/̖]0������9��uD;��Q�^���܈��X����	 -3H�����y'�r~�S9�]�I��g�'7n��Y�wV�p~���ؓT���\�Y���sd�51�v��=+�x=���<�����j�2�v��Xz^�U���
�W�@�-,�X��\�83`����Y���s$�\�� RV l�&Pw��>B�������,�n�����u�ù�s���3	�F9,��m�@��X �й�g
�']&N�-#_�Y�_C4�w�'X�h����� �k
w�U'�YpOKt~��|�l��:�����K�6��h�㚉���<�������q�ٍ����)���dU ����{/�U}�j�7�NW�?�L����������	g;�������i��	]�-Kf,��a�á��	gFѥ <6�Z�f�*�W��$�bV�j�`R~�:���V$�H�K^�������V�j���.�;֪�@�Av��Xle�?8ʀ�#S��ֲ."���[�� 9t��d�IW��RG�㧢me(Ғ�Z�l��`�/�牖�E�F�/u��3(-��朗D��ZC�[�q�&k��Dg���|Z�v4(:�+������=��{�N�sq*���E��Y�x���Ks��]�����<�9���X�e���V��b�L�ا��!��F�c�gi8'L�l�T�:b/��7��5!�������‒��hZ 8��ܩ�~��ͻ=�t�F��R72�v˔�؆������Qۮ��]�l��^6>,��M����޾魞 <]�5'6�
[���{��
YS��s{r��U�6�:��`�Krޭ��N�ځ��Lis��m�?�3����9�d��C�/�6;C���l��'�d�s�Ό)@�*c�{�����c�$��ϰx�`���fy$�K� 7���!��N5
&Nq�2�!�v��V�G�E�����z+�EG����X���/�5��KG�R��5�}�]Q]S/!�E�`�L	�4]2*�5���oBhdb�C��(؈_kG�^?(������s����Pq����Ew]��J���S`�V�9��3��+j��^<�/� ���ٻ&���Ç�ꝋTW����|�7�׏��W����ڱ�2�`^�����XKxz����~�Б��|�Mo��tOw���"9E�� �y@,lߦ���  ���;�W���H^�`�7Cw�^��N��Pd�W�tV������y�J��P��d�*�^b��;��QK	��ӗt�?�^W�V�@~��*T�/g
�Vŝ���,�.U���%��d\~����ZFu�3��/½ ���`��$n��l�� >�;���6l�8�R3$g���|N�I@U����=)hXqf'Gt��m�F�6I\��6I���� odO���K�!��������4,\����wߜ��+-Q����a�����I�O j�����u]o{�਄-qTWW�L��+
��CU�Zcޕ��w�����~���	�;_����x�,U� 	Y�ܔ]`���@q�ZЌ�CӼ�#X8����G��ösg��=����<����,pt�TI�)#$){��v�QRȗ��Py|����kMb/"��?�����C���O��H�0��^[aRӰ�*ݦ��H����k�g�llٲr?�/D��Oc,/�Ʋ�<�m�����:l�~�՞��ޕ��ж)��C�> dd�o�mm☚�ɩ !X3Eo�+�l�S����!C�-ղNӇx�P�����|�Q6�E����Q�r�x�e��O�LT�-%��Z<�/�!7�Y��9�)�K�KrɌ�����"��-������chR�����C0��U��y�xvaۂJg�����p.��	��8i�G�E�C]��L�$l���B�R�7�lH���z�NQ:�͇�x{[ͯ��m�2�@=Q��V�h����2��SG��7�A����&܂C�C��h�ES�Y�tρٲ,�0��NE�> >F4�>�#�-�sG�Ȍ�n�X�3k�M�.#{���G\W�z�:Ð�B�T�?@��蟨O���|�Y7�I���юޖ19*D)?>�賧'g�����L�U��v}�W�Pz��55��P�Ҳ^��5������c^F�j�ly}vW_�D"--�w�I[�9.�{Ar�w�F
C71�W��':j��x�(e����[�A�J���B��rjM�X|�E�z�x/N�vб��VIa^�(jj�̯���P����
Lg���VI��_G��J��r@��gԨ�`���3�Rv!<e�ld��Z���� J"Nę<��hz�C�e��3tC���:���KJ��[��ȇ�_C�l���n���.}[�~�l�1�l�ʪ���S���%��)���\���<��n^��T�������P3]e�%�!I�����?c�֗�@@$~���3-�q�}ϳ��%U��f��3�2�tA�	�`��zڝ:BXw͈P�̀�~�^u{�nެ_�A���q�MXt��z^`����9���N�����GCӭ4S�,	��»YK����~5��A��{��:�Z����&GV0n��2�Ʃ���~K�y\�������ґ����3ֲ�?�/�w�1&v*�ٵ����Dl�9�m,b/'�dQ��ܻ�%��2��ŐW둹�}DFU���t�B2q���D�|��E��)}��dp�
�ı�d$0���w���	����	����{��E3��o���_N�aW���z��}���m�%L�}>J��|�}x���?���9~~f��\H9�?�3�����׬��1����+��VϽʰl��Ћ�=
=����=������k�-��	�Y'hG>;ԏ��e{Ij/δ����'G9ȶw,�0���M����L��Bc��D�#�°�L@��@�I�s��F$	F�W%��1�S�9�@<���W=/h�X��Ե�,�"�>�8��qլj�� t��h�H�����X^$�����Ҽ�̽~�PMv����y�W9�_|ܩp��D�h��C�G8��5S{!ƭ �`.3e��4������_��]!]�Y�tgtpX;z��m�^���Xn]�\��hw�Ws���g���|�Pu/���B������rfq�Օfn~e�ތ8�Z�)S,�K�5��m�b�DO�l-$��S�Ц����з���0���%Y/���P����9�Y+{��x=1á�S��O�Qۛ��MM��h��G�n)H�����6���I,��,'-�f�:C�V]��F5��zDs7����A��L���k��
�՚j������$E��i{��t$��໌��@@D���>�P.ӊg� :^! �;,Մm�T4s'�����y�����muѭ�jD��T-�lm�dVt�;�Tu(�ݬl����H�ݎK�n�����ڜYӵ���h�@�Ķ�1NĤ� �"Km��1n��(�
��>�yR���F�IH?Z�¹9�l9�֠y���k�I�sy4NG�h����퀳��۟)�[[AfEp��$����EnsK���w��f$͖ռգ0�4��Z��Xcr��y
�Ot���ĦM��o�J%�m�}M���[�����+O�r�Da�����,$�#�s�{r��}d>%�|���; I�/����7�fYt�uj��X�t)U*3��t��߬�ܹV�|x����#6�@��E��Q���8)Fv-�ݟ&�xSj�T�*���4���TB��"�?�)S.Vͫ�{W��HU��-�tk���՞��6�T0z����[\5�(���hd ��Q=��x����/�im��Ȗ�t;)+Ċ�O�q`�g29���o�_k�	ߋq2��u����$��12"�o�R�@���Ncmi�����W*�z��6K�����l��>y�[��m�����F�h�\����&�PR����0V���Վ�e �P�a�e5����wHp��΁!��ǼV�������a�W0e4�pΔsC
Ӛ�}��҄���0����H��p�+�?��!L����1��P=>�6V���Vt]���t�Q�m�s'�{��E��;[��;S�֌_��]��8%y�⛆y���K�#v�������l�k�]w�d��vx�&��E���Z����k ��N�ڕ}o��#C�Wbj$qK�E"|�XDڮ�n�1�� aY�8uc�~��MU'v��:���-�/�J��s���>�O�,���"�0�܎w
]'_��a+"N��	�c����9�['-�ο��7]�j��ܚ�٠l�W����z'�6�Y���>c!��>lv�8B���ozD�0��`86�#����ƽ�[;�Īܽ-��$q�2z�oٹ-�N	�Sp΢{�Ls�$�����{#ʷDÀ���e]Y�X��yi�/9��J�S�z��P���
������r��D�l�~�M����7�^�T��/�jM�n
&���/�,�I�H`�b�������U�mC8�f��;�*��>R��:��	�Qzd~���u��*���s������Y!p�}D�2m~Sa;3P�l����������ψ���w��'�!QKZ�#l%���0�V�+�{(��(5B��Mᅔ��Q{�R٭�C��i�q�i�Ls�pK?��l։��֚�\����֡� ��4ߩ�����{I{Yb,�_�\��K?���>������f�eQ睸�1e��ɫ�I�����֎��k6h X6���u�A'C�O�em`x�q��q0���{ �K)q\-���]�=u*��Z��6�H�{�a6�e5�D.ä�����Z�X�aS^���A@u��D��$M1���T5��z�1�l+gPaF�R��=��g+��qV�ۙ��8��,C���":�a_��U:�׌ji�����x��U����$tH�&j��#I�~rńnrET��c(Q�}i�����j���˃.�z`�f6��a�D�}�b)�ô�\�`�`�U�^հA�T�<�+���d�ӄۺ� X]i��;�l]����LʀK��b�ܡ��ֵ=)���!^u[u_���9��cz��gފ��f����G�^܇��7�������O^Dݙ ����,�ޟ�цSK��k�ٷ���ѿ瑎"A#��MS|ѠC@�/�N-�(��ȱ���WRܼi~Jfp�ORwyHצ'jЁW���]%|���-��$��5�6r��I\��j�M�������mA%��k��4�V&v���Ӯ1���,�K�ǐf	�};od�ٲ�ߛ�(]�g`Y�ctC.��V�z%�fK�UJI�LP<�}��e55�Wv�7�6ӇHtv�q���q�^�"w��t�ڑo������VH�$eWÓ!���@��k�uY��ˏG����%#:
npEokCPk�'~CT�%h:�ۍ��L�b=�����4r.��G�K��.�����N�>�3�=���J X�̰��sܻ�}��a"Tz�b�k�
�i���R1ݒ���[<x�~yk���|�&\}��9n����k��=����R�X-�hЭ Eӳ���H�Xm�;l����7h�)\�A����>��-[���@l~x���Q	0���=!1bQ}l��y�<ߨg/���@��ι�=9��"������9�o����{'�o�X��9��8~���o�}q���bM�bX�x>}�LR�~�~�i�Ͼh�?�w�Ct��`�ּ�w�7>���p[��y���ӧ�`���0a��K窲�߁#tc��5.9ګgx
@�(�Tg�Vs��e�mV�dq�Bf>�_�1w�9��:�}O�7�f��"T�����\a!�?��0E�ғ.s:�yH�����]0�Ə&�Ox�'�!Z���9�ׯ��5�+��s�p?������)A����F�	�ے]y��lk2ӈ�vT2�Ft�#񈓾��o�f�� T��f�<�0���XQ��~��9���|�V�a	(8OS������d��K��	�7+-Ǝ�_�z�Ó15>�M.��l�4���&
�����p%xu=�,m�?�r����"���<ZRb�*9yC�42�??����?��������H�-�����uw;@��З��RY0� �&�*����X���yh��[=<�*�D�����Z���)ݹ�H�s��0;����!X
*v=	�26[7}�e(�M��MޏV����$GR6�H��1��*�h��a�;;���<kI��X3��؊@�S`��l ��ލ�nh��`-��H| L���^P�
�|K���{�=[���j��l$����]K_����4ȼ��z��~�:٠�唸Z��F�}���W��~�Sz/?�uc�������x2c?[���i��������r�5e��ȧ��q�}W�<nW��*���B�Oۤ� P�o��,�&8�	?iV��S����>�?tN<�u���~�	z������=?a*��U�)!���x���#O`
�Z�	K�#��K�n�����K�B��x�6�.�,�y9�k-pA�YJI�0�*�a�bM��^
�M���������P�NZ�+y0�b����4���e��'ϋ'�8�}	��ׁ�����W�!Z�,`�;�G��&z�O?���|��iZB}��*P%�
a`���-�W���R�/�9r3�_6g�\�����v�N���|��}R����]����]���^�~a~��.�%@�p)�Iҽ*��fYy�P�����+M�ܺ�LkI�ء�H����߂���c6��~�G�n��qH�KG��o�'5�����]�.)/�_������nn�Z6��ۺ'ymp�Eٍ[��4�2�K������W��~�,��33+UB<wȵn��wD�2���Z�ڼ�J ��Ǭ��r3<S��l�<����R䧙�<����8w6���.kM�[B.��cѵ�&@j���MB[�>L?I3gm"��fyq�f���pAbb��ƅ~x���nUf2�������)�� X]��pC��3�8\%�.G�\9tT)�}�u��8���!�'��S�[\'g���v��M\����&�)Fq��&�%LU��B�
^�l�N�J-!">9D؂���`���Z��pR� ����rǒM�/p�-�/�'�?f���q���NW92Ce;$�x�����[^�s���b��h���D�q:�J���r6�rxǾl�É�=�"��5��r�7�/?Oד���f�t\`��2.�q�qW[�;��񌊼���etm��Á��~j���$���Nd�$�bҗ*�R�`�P��H}��B~�2�q��6Ύ��T�qNq募���' ���J��9��T`{c4����dT��TxR,l�N��I� ��4���>�^^ߖR�����7�b�W1z:km�#��:q���]�������o�dV�o�L٭�?7y=�L�v��T�a5п���e�08�EWm���%@#��?lx�p���N;���us���0q/��E�*v��E#��%��M�p����ߨ�Y�ƾ~�O�6��`$�Ѫ�~d/��R�����nk܏/�F��|�?Y���?㪡6�����!G�sč\ 1ugF��ŷ�:t��9�L�)'��� ����zӅ�k�<��1Pq�KO���J~���Of���4�������I3u!\����J���{~�h�G��xt��m���k��ϕ��8|ym�#�GH�:CH$��5P}�r�f0������$���R3O礜�_Y)}���R���(Ϫ|�'�G4����͈mn ^���`�W!��=�=t)�j�^Ģ�11�x����G�YD㣵+�=�zT�z��Hlߪ\�hFb��.}��	����\�[N�]��M�<\a�2�����c��7���������ہ�*����m�*�>���n�Ts����@�R��->��x�Sql��m�/� O���������jI2��a���?�ѱ�'�HǦ�Q@�����l�RS�OW��l=�7o<��c��'�<%�j��:��|�� ?��C-t|:���h�o4s�9Z῝����[Y<[,�^!��H��lUH@��&���'��%%R8]�HJ�]ۿi�;��偀^�!K;��[`G�~L�f2s �&0�Gm�Hh%�5�v��Er�=sS���.����[�zNw��UN�ě�-���4��џo/e��@��zD����ZF�X~��aN埍dO�^M?�ٍ�=&v؟r�a[����e?�+�{5��� -n6�.� ���@-}?���/v�J��~$��j��R�\a��/xWE �z�#�])�ص����G33���Y��@���{�J�P*.ak�
H�}��1�=�f�>xt���R~|�m���q��W1�QzM�x��;eLRH�ҟ�E���m9˒��aA��@��##�O��Հ����b�Ҏ���2�zL����G���/�^�3.��_udJ���t��/��nA�����X	���:1#N��{Pב��O�O�AMu'|f�=����Ͼmc�|đ�,o����X��-H���e�AB>դشR���a��SUr�BrxSj~K6p��%䚑j��:���RyZ��fd��W-�AW�;ܩ�5?��C��!Q=�x9�i�Zi�W�jN���v_K���P�*�)E�w����?�o�%O/!�ܗ�7�ædD�ɗ���W&w�_m����R����s��`��7�o+�H���"X�2�?�Kf�&6us{q�����R!�xv%b99ӰU����-J8��M�|�� 7�H��l:�:������=O��]P��QAk�l�����܂��&���|��S\-y������}�M餗��!�GL����HCT� ]�0̎��;��.^�ְg)�l-�;;+�wF����q���*�����`ƣ5�@�k˖���̱��"s���x�|e�i����&.R�We���깢��T�~��Dl�n�ې?�3�v����Tr�.��\����k[�2���(X���I?U�}�p�W�Oߌ���E����r|y�ef�J��մ1v���i{mq%��֚�YWMl~�B�[�p;,o�Xq�x�r���`�׺6��G�&�8¶<ܙ��@� Z��'������$T�e����f�M����_"LP}!�U|IAU���B\����v%�Ba���>|�x2�j�%�YLL,1��"l_J(V�Ʃ���aȆ^�<{��"rul�Z�}u�m���s>5��Ń��˹8V����rW*L���0G��8E��)�B��A��fw~S�d�S���4�- 3���X�CC�I0�)ܽS��?�z{e�&>��
�l�֐2k6�W�����j��h�c)η�>����3à��T2!�M��e�{�ڛB�YŘ�+�����sv}��eʍ�7v�k��{EwV�6q!p��O��*��U��@iC=����� e�5��]U���N/l��is='���'O�É��7��+�E�󎤜)g���z=�\y|�),�;udSа��C���Jf�>�K��|��y������#�C`��?�W��YN���Lt�D&���Dk� �z�4lR�W9-�S�������2=M�kSt�43����,��#�y� V�_��[��} �8r�l�X'�{]\+�~im�>I�j�wt��5��,���g����V��h�>1�*�2�g�/����i࿵�/	���
��#��D�j@	��x-WД��ܠ�K��kKC{{]�4��F�)|:<