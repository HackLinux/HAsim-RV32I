�Q��)a^01����
!)�j�(	E�oJ���I�,6$�y��t'2��\�D��<�&��<�[�*����2e_�@��%�9D�R1O���A�Gu$#����c�H'M�}������*F�(V?i@V#���\��kL	�>���OV#�5 NRZ��:H'sE�P4)p~ңX�4&��O&Լ�����v���U����d�<��V��wPI$;�0Rΰ9S�/ED�PDF؜��&9�$�i%���!�Tz��A$�7�(o�HAU����^vY��L�G�U��bg\�-�����2k�'�[��$͝�v�����NP_t��ؖ��\aCfig��m�֞�y�,����X%K;&ӍĐl�$�0�KK������?\�%�cu��wG�$y�]�oO�B�gi�/b�k��̿8w�эAL7��;"�ӗ�tA���r�����j�P"Kq���E��`0��n�e� �%��o#���hNAW.e�	-��?z�w ���d�)y1��2pX( ��2���L�H��F���F��@���%)23�h.S�����*:a�DFMǏVpd\��Q��l���p�2ia-g��%E����?�FٴUƠ	s�Ҕ���e��]��x���j��I�y!Q"s��3��A��<F�i���foPF�EGX�?+�L{)�����5l�"w�i�� �h�;�6�r��w��UN�!^"W����Ch��#�����H�ov<ĕ^�`�1NB��̒{����p�svB�� '�󒜱͜0漂�t��kd��0/\␊<�>A���d��*]��Ԅ�g�C0�EuHpa�dF�b��a�r��*U�3�7H����4Zx�VvY�]�`��w��������Z��T�B1?�Nj���q�/R�!$2.�Z�
�.*�OKήb��/��jNg�h�#MY�Ir��lb<�-g��ks��!��/��J�]��m�jH�2�F�1:u|S���`K �-����K�R8���l�ECY�o�HUG�v* A�g��u�i���_*{�Rk,����@m�M�[qSy��pO��@J��ܹ�9�a}��V�/�S�1\.Ѳqє��U�rƨ�3�	��!fN�	䎝0*j{��A��C���Iz9��v�ڑ�cx�0������87_k[��!��A���ei��ԑ�.�Y͠�7#�a[�@[θ��|.C~���C$Puw�/j�A7�kI�J���)&�P�"~�8��䙒90<d'Uy�*Im��V�-�rF)�U�@�m�m�n0�'��E�*��MH-�\A��">�o�ʁ����i���#�bb{u2Y�ΐ0�"���JR����&"x�H�?�֞�&X!�4z�4S6�j2�WN����8r�jڇ�+�9�B
a�e� Gˎ����d=��0�����d�U>*5A��,�4$��8?E��΋�琌8T�bQ&,{5A�>BY�p��\�I�y��Vk�,�s�.,D���&L�kS?+��"����E3,Ƨ�:!uy�ֆ���%�����i� a8�oB�l��"�p�)I!v��}�.�Q(��u���vK'��M�8Dl}ks�Gc4_�̈́G�
5K�"F�&������T+�ѓrQ�c�D�U�OGp���3A���+�xBt�7 �k�����*[&�F1���U�aAH"(6�H��b��Q�a5Ҫ�����(g!�DVͳ	@��یV�w�	�w&,�o�X:��r98�xuע��,[1�X֥a8��Q��5LP"�0�M3!���f�ci{��F�אwUl_���E��(໛��r���-Fz�C(���䗬�2��r��S�S{U�^�6ԑ�Q�jH���SJ"7��i�$:NH�Nq��H<�BE�I�JÙ��Y��L#3���X^��)3��X�8f��YK�������aVfdV�4dťmk��U��圜Z���3�O[c4��̥\0x�,iR&�'�?�&�L,��p
���p:�N�K�,��)�B:#�-[�t�4�%K�b�h�L@e��2p�:��%�@8����SK��<)ҟ�ұ!wg9�>���\��o�LnS�Z�!R�D�tV,�#sm�T
]+�� ����=z�V2Q��R��t�t�'Z��꣦JSJL��G�GT$b��2�iŤ�^���kEw�⻷������;(��cV9`�2�B���,8^��Ve����� L��bIju���|f�6@fb�U��U�%{5Ȳ���*p�vn�j`��]U�\�$����� ���:8��]�Z����ո9�J��@M\�)=鬔`:Օ"ge���.�K�K�"mF���Bi��fil�!Ҳ�X�=T���s)��A�/��u�֖0�ەݪu �%D��\4M�����O阓��y�%���I���ER����f6��e�.G�f� :�)��8\[.3Q�����cV��<k�1Gol[����ߙ(�����(H�/]Lf�F��O��71�Eه�}��U$��z�������:v���b��l��eÝ�A�3�eH�(���f�-���2��m�@nT�N/���g\ƾ��6_�n�a�<���$�9H���s�+�/�̗�(,��}狐���D�:;���B~'�:�D*���*=X8�J�*�R�xGe��g�ep��w$��I_�qTj���,�tp�W�[�|+DTM㴈\�g��ILjŎ(� ��x�g"�r즪�H��HW���y�Ȍ$�\�\�Ų(�c�1rJz���	*�s|C9�A��\��X���BT�s�켴 �yt��Htw����&U._�"�p͚IK�E��0mA���%C�Љ*dG�C�~�t��uǈ��Gb�@?��>oԏܸ7��@O�ӀF�Bdd���-^d��#%kE�"�&+�VB��^9ZGdO��Q���]����)Nr�i�dk��IV�E~�YI�������5+煩2��,Z�%��#d��l9B2˽iؼ�nWYܲ	�!9�d�-����#���e��F݂���[��\}9#�HxnHAt�f'l�	g�OO �|��8Ē��R.l3�(�-�	V��5i~��*}��ΖO�Y���0���V��jZ��e˱jf^y��c^߆���q��[�hTo�
c�H|��y���2b�v#�+�R����)�c���k&��4Md��tAW	��rۋk��nlZ��(�4��9�
�Qpl=�d!JBc�t�:�:K;1owЯ��y�ʰ9�`xca�����8�lS7�R<�T��hc"z�b�1�]�2���Бؠ7h�<U:��2)[pȝ~)��̑�̼A+�}��/,@N$ �8�D[�I���
Kr^�� ���tB ��&����P�m�,�Z�FR��7������g��)�|�gK��q���[|��H������G5�Ճ)�-F@`���\͖Z���@ 6���'���I� s��^)D"��e���{5�hA�"�T@W={�N���m<D����Bk[.%a�inK!��w�H��`�L��M ��H�QƱG�<r�+SK�;��6�"�د_��7F�!�[���_��VV<�ݩ���N�~X6��68�O"��`��Th1�E-��D\Zc���~�9bY�8> �1y_��U�յ����wK��g���<֬�T���JB�$�Β��`�X�:-�uU�[;�;ۻ�W�� Ry�կ6٫�Z�l6��m^ֹz��N3h����y�k�pۨ��c�^nm�]������e]���J��V,�xyqms�)�ܒow4�0�\.rRDLD�b�j[3 U��Z����𾔵0*�*
�p`KNpΨ�|<�
�$���К��R�ıSq�Z����M��!��'�k�`������Kii���Y4X[�B�.��Fj%8��0^�iǜ�%������p��Ҽ����7o�Gh���R�C�	S�E��i��z��)=}���4&R�� J���8
� ��F���M:�o�0r	b4o�t4��_�pź��	+m���2��jɢ��$�R����+����JT��b��ƒfg��78�?C8o���{5��X��d������9���o_���̚�%Ǌ�\�l���B��/2pX"�ɿ�Ҷ-����+ޡ�B�q��ㆱ�b{�w�l3��UBr��D�ַ0k���0���E��Y�L�|m\:����{�K9�0����[��|�+�8���:g������mnq�9��#1�k��^Η�V�XY[l��x�1���׵T4jc��ڥ�X1�h/�^�R�^�xEez��V�.���a��_��4�%F��+�i�"�RP�괞Qիh��B�9��I
EM���:�����h��x9�q&^<~� ���pZ��!���b+�����-9�˅����������:WY���OY�l��ˇO!#��=f��tj���R	��˪�,]Uqx���+C��]@!�IKu'5�&v���i�o F�y�IX�xn崊����{�f9���6�cky�4�֯��]u
���k庪{�б�s�d(�o�X���u�0�Jv@�:��R��f��9BJ�C[E���G�A�akd9���t�SK����#
#M�*`:A���D��g}��76��4�`�j�<?��p��9wts|9�p�4F�h���ȑ�Xh`��ʬ���jX��ְ�4ϡ.��8}�!RU[̤dV�LJ���ĥ���r��b}����˲�^��X�2�CJ?����iͺiP�ҿ�j�no8�o/��k� �\Ѩ�Q�V>��1�������0���U�ZtO�ҥF,���>��$���u�ǲJ�K���b��@Vj�l��PY�����B��=�ֻR�Hu�(���9i+��U��NBD(C�_q'�M%��.��LyRU�t�]E�+%���u�#A�1��IB=�©��td�S��c��*��t��Q��