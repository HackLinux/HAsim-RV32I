�4`'�����:oOJ#��$�	���I �N�W���O��o@��)������d/L�b�g��t5��E���umF�W$�q<����1I�{6��Y����� Mf�MI~�?܃���N�a���.�O���K8-F�������3��Y�<n��EȎ/��>�B�wݜ�a������m��
�≛5�/[ᯆ#�e�,z�+i�y3������g��]sA��ҟ�o�AN~�������3>�_�E2��L�f����D��� �/|=���Q~�������H.}��S�''��a���+�J�]a[�%9�{s�i�ۿN,S��q^�Jo.K�#�皤��߶���/#��=n�=v�]�C7~�?�n�X��ek���$�RR�Q-������`I./�M���g�y;wumb�\}���_�����3=���o��]���&{����W�9�\��^�a�6!q�K��*��-��`���0u�Y��_��l9�=����a��}5�H�%�iI&�H塛��������O����#��G6(aL��T��N�FjB;U��p�P�˾lo*#d�l=#�2��w�?}n�{��ɟ�sy\�-����(g��f�FKlĢf��)ֱ]_ķ���b�b|z7�s�E`Z�;��'��J�c���3㱾�\��o�KCH��Q�!��*N�=ǿ��Zu-G��[,/�8L��]�"�����_b�����n��O�K���ƭ]�!s�+����~R6~�k�s%|�9j��5Z���tY�_2'-���fDk'��u����9�����ϭw����<m>�=難!u�ػ�����Zi��$����vfӂ}�e� M߄V��'8�(YS��؉Gy��9��ڛv����S�rp��F�d6�8�Z!���
#�|��g�[��9�L��-F4Ç��x~9����~����וe6/�ԗL"�� ��5��ε�m�b�>����Mk�%�i��4rf�2��UW&��<G$��L��螔>�!,��c
8�iI5Dw���髾:�hZ�M(�����p��RA�ǿ�6!��ϧx?r%?ھ�8�&{Ty�V�CN� _�/WR���h��sD��t��5�i)p���I)�Wu��x�n�΂���a���z���"�:N�d�sJ�k^��em��;����M���J��m[���Q2�q֊��9���D���/_YVz?\�z����w�v�>Rk�a����]���w������*ĵj��=7 B��7�:m�Q��߇�� �n������k�=��$ �v���5�JXY�5��8B~z��sKD�E������T�Z��k��g�P��u�u�?S)r����95�yH�Q��}�FL|��z��u�H\�P��u��x�i�\nݧ��Gh�"��߯�Td}��Ƙ� ��(�E������|�,6�:a�g�����j����~N����cЈ���v;���
�D�Ȼd=�@����j�њ�d� �TW
m%�=���¡r�p���P�1��QR�����<�!%�4�;\O����?��Z��8�u��E��%_���3ᐗ�S�������7Nk�OSDW{�79����H��%3]kn���~�}|(�א�vl&�����
�*_CG��/w���Jo��èQщ�����V�mC$uOH���}Ѡ�������
qq&��5_�:i���O����g��rK)���B!?�>�|~�nV�}��F<!��o��R��d|挠�hH�?�)�3�~x�v&pߒ{"�~��=~a�e���S��y]��pQH��Q�t/c�����I#��.�aԌ>�}�s���y�I_a-�^��-����_�Ng]�R���юM�vWoN�6�cR�i ���Z���L��} �V�q.�z��J���[i-V۬
�0��GZ-�E���eCJZ��ݵX�~$��IѯB��Ny��V�h�R���n��D�E6�>"k��Hdɐ3�Go{����0��ͪS>�`KICֵA�S�q�<�LR���ؚr·�o��=C�iY�1U��e�W4 9��i�ϭ�f�M�z�}����'<�D��J.����A%�R5�C�|����/�v���h��W�J�,�[D�����Q$��)#��p�ߊ;�]�Z_�A�^N
��k~��\n��F�qK��Bx�����^}C�!Zڡ��LW%�&����;�����ذ������ 22��c���/4'dNc�����Y�c���G�]�� R4���&BI��J�b�ݓ|���b�#MI�'i��c�� .�"�M׳��7�hҗ�ڋM�S������{�d��5�i���-e13|m6�%��9ԆP:'
��F>�V�*��:C��j�~1Ȑ�t�bh�d\���砽��S�d�u�~�:%nf�	�� M_��I�Щ�,Y\��'`p�&���g�y3RT@FCՂ ���GyG�����.�&KZ�#����U��v ��B������7�9��{59���.�e��;����N7N�y�����,���78�f�k(vH��H��-G���8�r�Ӥ�N����C�3�:Q{=�2�:�����������{�)�1g3��N%��ߜ��a��O�>7��J�����L��T��?�cs��zz~���p+{ο���O�����zE+��Zqf#�fe�}���^_3�wႌ��R��x`���s侎{�g$�;���
�W��3��J�D�愈�u�3��|��1}�x�)�7�iE���I]j7?E��jwN{X����É/XGo�3*FX�Oj� w$c�,��l�֚+V��?���&����q�=�&�>'Ѷ�U㷆g��am�u��iH+���B2���U0C{��5�>ŷ�V���Ze��p�.��i�ۺJ��W�K�毣��G�a���ƨ�H�L3y��K �lz���箑+Y{�� K+q������@m��+���/T�Y�j�о%���;MSt�ھx4=��9w����9�|i�x�H���.� �+���槛�bX8r7{��Bф��(t��ݕ0��;LK��]�����S��>굨��{¿|�a���"^@[�8�Pv�G���O_�?����M��7���q��`�]�N� ��x[u0��o�*eC�jʹ��^�����MZ> �}�}�җZ�@ɤ���h�0t?��� �Y�Q�ҳ�77K�T���6���׽U�a���H�R��4�-�z��|}-x�:Ұ��VY)	�J�Eǥ}���U�����e�g�{Yݣ�X�AЇbd3ɜ�іE�rZ��G�tx��^S/�/�?���H�������ʟ�:�3G�%�3�%�[�
�#�ع'��ǥ )�M���Qw!�%��BZgy{YTp�x��]�Xݵ��������Ѕ-od����ɼ	��T��#}��A�e�������H�4!���W��*�8F.}��Y�k�A��[�/�٠&�4��~�iP�*�(�0���.��-���`��K�OU]�w�E8]���!ggǿ` �7�LG���h�ln��B���/c'Q}���a���ī�51�����`/J�O���:��ew�������eZQ$���v�o�*������006��$�ye��+�<d�O��+�a�-������:��;��H��M�d�,ۛ4�+�'	��}|[�د[�g��oCL�:��C�����f�o��y*��.����j_(��g��W��wޢo���wQ���N���t��O�
�^�Ŵb5�֛�^�y�%-�%/Lt'�:3#w�}��P�%��/[���B���
����dy��&�"C��d杸����G?��T�Cڟ���^���ͯ;A���y-܇~����"�U���b��>�4>22֨��;��*c�ڶϼ�O�Mj���5����&5�����V���a�޵Nwv��䚠��R��%��:7��یL��7��#�K�ks@y�����p���4��uB@� _�B1>x{a��,�
��d�4�E�j>&u�&UQ��Df�o�D=��f�_��@Y� ����y�;�����������_��G���7�1+�>;�[# �aCX'߻��������U�����T#���j���p2��1ѫ�dyl)5��Lh̜A�++W09�k�
7sz�0%�p3�W��t���R'?�E�í�W����ʿ@��	��-Smj^[%�MP;�Z	8"~U'&%�M'��=��豴o���YIw���=���τ��J-�����Ex�~V�R��}�Mi�A-�&	�/ݚ���Ci8Ǘ�L�yCP��I�i���i?�P�T���Y��1����x�N �a{��J7;S�
[,a.<�ߤ�y�1z�"�RN�d���C��4s�3au{$�W-S�j.�[/����q�M�Ș/l�Z�������vaVv��u�#|�v�,�YkDl�ô���m����5���
K��]��T¹�m�����wg��p�=xU2#�sʯ�<�Ɵ�xb㑕�����w:��cp�@���>#_>�φ�xwbzJ(_G,=���OK����d,Z�����z��&$���ȹ�a7]=�]�"�umKQwgb1j}��T�e�s�ߡ\��ا坿^|�dhi����j��56_���&�+q���O�0��2CiE�}ͱC4�z;�#���_Ҡī��D8�+=�,����i�����?�Hs����%^.�����C5DXZ>��d3��X&o��y��9�)��hl���H���zao�jA�D GQ�52�	�o�ԭEE����~"��~��G�0��������;��4g��H��o�9H9'�|� �QvI�1&(�C�R�����-[�d?^f��^�u�_*y=Mww�{ĝ���M�N�Y�`t�X� �L���4�ִ]� �����9"�(4Ȣ �S d�}��A�D �<]��L~�X�*+�o��L��KxB_�}���d��[������$?#���ou��e��m&鑆a��>�Et�1|��	���rF%=�]�]%�������6ħ%Rޟ1�C|Za;l���ԢH��?�r���5ɑ5V���AYhOeX%��9�8S&8�m=,�<���-������U��*�<Tҋ��}��\b3�X�+R�=V玭��s�r��m�tw])��m�>�g����=��{/��c�Fv>N9ڞ��ߓ���uv��Ϥ߳%��.����l��c{��v�\h{����~�oy������V��a]��>�<�:k6�s�6���LC�)�V)�/̕��_<F�E@��=F{jM[�
���T'����B1bd��f�������kd��N ��
���9�'���ȗa�$�pOQ��,n�Y��C�̰��Pf��\�EUX�f��}�2����F|8c22YY��@�B�+CHe����u��Y�2+�B\�(��K$�ݤ~	�,n��5;aU�,n�4,�JЦ7�ˁ�z����ea�ո�'Y�H�E��Twa�x|��]�C³�9�n.�F<g��"��-�y�W�<��j��q��#o�ƃ խ��pK67��!tT�0F#��={�.}�Ɵёn�0���z�;�ş�`Z?C�!��某_7�)xa�ТEG}x66�E!�Tz,�� �nO���FH	�R��g��3]ō�A�������C*���`z��Ĳ�m鍍���@�TE��EOHu9t�jhTS�X��޼�����}�e�r7�@�X�FeA[��]���&�m
,�cwj;�XB��v�&�tv�2��-.bۜ�z8N�Іa7ǳJ	?�
��=1ǫG
,���0�2�Q�����W�М��ϸ�t�@��}���=��CK.;N,��tO���F�����(��U�$�~�Ph@@d��׎�΀�.,%'ڸ0���s�h���=](E�ҭ�x��
,�
nl�7A�=�Q y	exF;����$�?������{��E���?�@&���D��~� �0�)�;����u.ĝG>$�+#�n����Ew�^G�� 0�_CHh��f�0bp���.B�!Z=��v�"z��T��U (�ݭ�]�>E+#Ұ�s�"$���|U�T {�>3E��d�������VW�����[��{����(.���u�6=�h��=Y���YV��+�(���jX{>5�t����;�����8�x� a��N �	2�y��s4���觡͌��F���UEY|76�>�X M�$\�V�j���V/��9p�k���+A��)�����p�5�c�*�Y��꜕1���X]����A�8ۧ�4����K�Ҩ}6���8����E��@I�0X��e�����-{4�~�t��:��G���*�дU	��}�?WM�s�j�X�H�*4��}\�\�� _ms���^�d����	����]��]��� {��$Ӱ�<Z&2 ,����VT���ݞk�x��{f$��֤��"�5~Q�UG��&��7�6G��'l�4�+4� ��9��-��C���"ʾԐM�8*�!�xm�>�8[n�r���@�]{��e�G�P;�l�����܉2eI�N�J n�sC۝C��p�¼H*LЕE��Ӑy�A�¸�۸V&CY� ����M�y�	�i�#Q�k#�&����룠�^:2��c?Z��uG�~X�4���o6oq���v:���Ö�������H�̈́�TZG k��Gk	r9�P�6��P�ݵ���������G�	!�_�u�$�T���5\�C}���0u�x�(}����� 6�d��~�5���R��X����0��������;9J6����A�(�L�)��+�31hR# ���v^a�e��I�mA-�`�)A�v���B
���%�-�����[%���g��7���G��Y�J�d@��s��z��y�t��<��j�^l;��1e��gE6ǽ�iK�yc��k�ό��h˚� [�BZJzJbK���>�,'G-��(޿`�i�ˣ��S �a�ja���sfTaxPVD�<�<�y�e���]����CO&�*�� ���:w�$�Z��e9���T{�0��dT|τ�Yf����oC��QWVgQ�"�󾔤"��6���D:�&쌌^�.g(���B{l�#��n�^5X�\r��Wva�]��(pE����I�������9��N�����q,���>�
�t�J�;{��)
�h��� ?���k�7��-dH�����a?�1��wK�\K�q{D�������j3�u4�q���o����Z1��{�u>�^E�,�p@9~z�|m�+��>�(�Ѩ҆�0Sc� �*(�O� ��6����M6��R�R��l��g���K1!K����uKB�yI�fAY��ۈ���?y��Zu��㏟�*tA����*9�)�P@�Z�F�0��75�Nڄ����u����І�s�v1jm�`rO�\�Y�\���x�p�XB�D���OOTN"M�'�$G%�%F$�"p#/"�#5"� I�v��>����?�O%�+�*�1�(n�"�<�Z�D;��L�L6�R�n3Nrʃ�R����R Ì��dT��=Sp�[��j�2�~	��QGڡQ�t�VN>�wp(vz�T����84�����I��xR{C�\�9=���U�I	`*��8�D����M�i�X(v�!Ӎ����h��YT�DD��e�� C�=��@� �]�(��֊���P��C`7��B��uD,�����Q�+����SZ�����k�}53��_֦4�Ɖ��/.��BNd�+3�p��8��WZ�K|�y�Ԇ�	�wQW���P���Ć��dY�(��7m��T�2�sN?�vx���Y�v=��@���4�@�G�@H9���ګ�#?-
�X��[��eU�d9�`PYΣt�ܸV�`�{�9��`Q���޽�#�v���������C�dxv6B/2�`X0vn�@�
���4�����$jPGH�'Pέ����P�E�u��������B��zҺb�9)#���������d�􄤥T�~
ZO]=^ |n@�B5�ת�'êk�ׇ A���_�?s�������w���+�����K��G�#�#= �|5|�o�����7���?l��,�?��/= �^
8�>�� �� K  �.��Ni�; ����|H����C *P	F -�iy_��B��o���Wv+	�2kO����1H�Z*w͝��^�� �|'����C�C�"����5ZW�Շ?^n���ҁ���7^�'��FN@������~�����b
��W0������)	��}�܃�c�$�9������o�?V�l�s�'��`�ӷ���@y�P2 /�I: ea]-�VA������D@�}L�|=����&��+��U��� v� �����n8�Rt{j�r?��nP�<�E@��po���n����"й9��FA�_�8w݈�-$�>��0`@ePtƩQg�Wn�dM��;�?}��U���?�r��^��縉)�!ϼ'��[ ư�2��jf�syj��"������c�q�
�K�O���:�4�ք����	�!�{�z>�g�i�^�ݛkI���-�W��n���#S�����B�9�Pr7)%P9�_Ė8����y,�.�RL�bZh>6;��F�-�Y��=��Q��!(�p@�4���������-�͓����"e�yh�ԅ��rs؅�K��h�"���w���R�-������T�>��B�Vm�-*N"g�W�ڪ�[��RDq������rϝ�A�eM׺`_g�;�j�ZN�S���lo��8TSD�e���a�+/�5�0�H�M2v�ͤ���CC�V�z;���g��j"S�uҐ��'ڏT���0<B��*W:>�����R�\ˁ�T��g��t�A+X�Y{s�%ݫF"���7����\��S�&�+���D�ἒ��0��\�j����q���Θ�����,ھMYB��� A�������!8+��d*��[-���郾Z^sQ�n���r�w|��7	Ṡ���[`Ҡ��w`��Z�HB�#nUvP�K��X�*1Un�p}���WL�7AW-�p>i��Bh�M�A1^l܀CX�X���ѻ�^¶B�]��yq�����s1bg�ht��l\�)�nc��<we�I�:�xvA��H��+d,�����	��#��� ���FO�@9Oo�Q���b�y~��x�^��;���;��`��ڟWᥲ��0N�˄��r��ϑ�L-�y��+S�ljj^<���������x���G���@��6<�%�y�nq�s�?b����a�d��/��cƢK��zM��K��eײ�,a-�_�i"�*��U1&��Qe;z,b`�~����u���E%��(鏭��[�2C���n���n�87��/���9߶�]��r9e�Ÿz��&������2�Y��_��r��F�cx������>Ѧ�v<�_�pl��B�� c��c Jc\�p�E���gd���L;v׻�DB�s
�oƫIw����i�'������6)A#˿���ĬC�?�0��G�6/�+g�닂x̽TS��u6]�r��<�~����OG�kQ�v��'�J3�L�� s^8F���ލ�[sX���ÚKwN��g����I�Wq�=M=�*%�!*AԾ��d��W6�EX����b���
�m�y�G+�b`����;��AM�h�gE�KҺ��ޞ�J.���w�?��etH�n����R����G�(��d�9���Y�Gf�w��,����m��f_<�{UȈ��a��("Jٌ�uxJ�����ʫ ?������bWc�#^�D	�����t�n!�Sa�K=�{vڽ� '�F�٢��Lܫm������?�h��{�9��h����b'|Mu"e^R^����_����FEBPz�|W^_��O�7�����l�^m����(N��m�AV��?��&ƱP��>�׺Fz��9s�e�56�}�|мпgzs��)<��G���&�"v+{Ze!.I�#r"e��%PXp�|*"�\<o5��2�KHteW��;o��x�g����>']V�|���C���SĹ��$JS�����xC�D
x�;���g��8���8������Q���M�U?��_wN��m���]�v!J���wu3oDA��a	�}8<?��o�ښ�/���}D�'�ǭ�{8����  �w�qȄ���n0}P������8
粂ۉ�M�-v�ٽ�B�_��U���u��]|�*,�� ^�n�Jy�5ka�b;��hJB)�1���G��M׋�e�@ ����]����p���/?o�yjq���9L��]�/,�I?�/՘�q𻊇��{P!�Y���8�'������k��7�;)�I᪋>�S2�B}�I�X|�ʚ��q����UD�(ye��9��^N����5�y{��ś���0�!����<�%�+M�3��:�z:���j\�X��������|U���q\�g��0�m}n��U�/�O"�
ϪW��tngɳ�˿�8��h볁U7���b��͛�q�̈́nh�^���sX��9�V~x���*"�/�ޥI��!��w0ȼ;�\���.p��'�����ۇp^�򱁌��1K��Uv��uʵߚ���;��XL�-�u>a��`�1�\v�q��xbf/ѫ��Dx,��}���F�r�:f�z�������~Vf����y��3j��u�ǐ�㟃�mYq���l�9�0)�$�O��!N�pu��I�?�9���#-�W¥�t��zl�9A�w�.w�˝�j�I=������u����28DU�
w�ܻun���'z���9-�쟖\��*­� _ZqH��^]��T�s 1�j�o����$8|���?Sz%bΥ�}�����alY��V�x�"=n��лk��~�\2�B=���z�_Fn5H��6&ӧKN��wt��q?%���|�x��p3ϡl7�4�=�}��.$h�ݧH;7-���������$?��a�y�3�������>y���b��?���$9���N#��廨O�(��+4J��a�]Qm�5��l�TcTC� ��8w�gZ���g�~P,L��A0��Kp4�A@Yj����]TB�L�d����:�~��	� 4��'���9,~g�?�>�{�����Ѻ��GKV�h�kOu���Q��������ؤ�&y�m��l=ٔ�/�����7�b�c��&��9yď�u��zⲂy/m7�7:x��f��ڛ/��O`*��y�VQ�b+c���QT��$"�m��z����p;���ݸ�n��4�:��q�����o�
�* N��I��k���"�!	�	��6@:���>i����}���N�c��-��{ Avg�V�|M���0�!O�a[	��$D�7���ꞧ8Q�"�6�<A6�C`�\u'��H#_��Z���[W�M�9 $�}��5��=,�A��b(	@ ��|� � 6��@�@s ��N���������\�.�U�7�K��� �	x�aM�-x�~�Mm�+8W������5�}���^k={�g��x�-3�<�7`߻�
��ͧc�5�\���k�ǹ	�k!ػ�gW�v%�n����7�����b_���eӳ���k��v�;�g�Xpn�	�\&���k�/k���^�������g��{��w�{���v��x�5����� ���� p���v�k�^.�şD&ޯ��g�[�_{m�2���� ��sr��|�͎t���~���LX�W�]�A�v@^ � � ���m��g�CO � � ̀� ��D!7�'}��F��~��o�����2����2}��m�`$~ɯ�׿��o��X5�P���l��)]S>�=�V����i90��Pۃ}TF����J�*J�Ûy�y��O��V�J���z��'K�@O>�XBl��<�f4f� ٚ��°�b7�{�7�H�� =^�X�>�ski%��|6�ʻSp8�ix�t.0ţ=��+6���
|@N�&X\�����l�Q��M��[2�Ȝ3��S� "���O�~UK��[�@V@X�uQ�Y��F��^����]qc�,� Ja?����z��~��p��q'�m�ݸoi��qW#wB�;���Q�*���nh�Օ�-����v>�����{��>{�<%��ߎ��UD� DT�>"D@>}�˝A��  A�p]�D}	�V�Q���\�D%� �����Te��������1�.=����2N^��z��%�G�SH����eb5#L�6���p/]Te�,1�dB�~��vKurY��������I����N��)IU�W�ͥV������t��D�S��4�2zR�1�%�VU��$s��܋	��d���R��{#P5N�X[Tƻd��&j��m�S�ty��LS�=Ljڵ��'�w�fF�`@rnk7��sİ��*�����ڕq���g�(��w���cE�jz�8{ĝ�l���zw+(��
���_�M��/�%$ټ�.�K���g������>VT��'��n�Vy7� *���� ��E��i`�/ X�x۹~����Xd�(E��9�
��:�ѻ�g��;3��` �-$Pp��y�����V��A������
�σ8Ab��z�(�+�0��	>�9�ӓ�z�xv ��J��Z���K{{���>f���">����I*˛��8����F+���߄��%]G��򿦦��$j����&����U�:�z0�
�<�H� ��'�tU
I�/,Eۊ~�H�ZM\x�|���R�Y9�a#a[�j�m'iu:5�f��!�y��N�oI�uXJq���c�U�?PMFm��c�=��_%��m�i:�>��z�)��p�����f��|w�ذ�m{��`�{�.����Gqt��׋��qS�4�ˎ�����z"�|Oܻjxh����c�L���Uh�������C s=�듬;���Q��9P�T�Q�x�i0���I�KFV@UUB/�{���?�.��tp�Sn�[�j=�U�
�����+�*�-��]����
:���.%��m�AR�u��q����ר�G	1I�}�w���������+xn�*����J~A�3oW�<�mq�U���<�yuȃ��#�R�����+���?r�2��
���9�$ї�A8�"��~��aȼ�����ߖ�漾K�?���(
	���%��T���J�+y����p�KF��d�6�G~Q�AY����W�v ŸEtnU��<��`�nl`�mis�ԩk�K��d�2�N?xsa�;���;��ހ�(�?B���7��uA��OM�}w�;-�g���\�]��]?)��D}����-��v��3<�� ��(fU�sl�� VO��g�!n�!�"��/$�;>��K�O��.Q*Tl�@yvv��O��y&)�v���
���@��͖`{z�I:�ů߫��V,��M�K�VO� �@9��~�H�� �p���'�"��� ,_;�Y�مH3Y]��ڃ�3�[��a��<QNe�<�Wh��f���B��F(��ft��ޘ^��S�W�a?�)G �~�D=i��O�Hə��mv��?��񌸖��|�p��C��W���}w�/i'}v��JrJ�����u:��]��Er+�p.Qa�0��k�n�o����<�k����R>�ܢ�oj��
�Q�{>x�x-�D���| �/6�"&�}D��3�o�"��2������)�zb������4S��g��wb ���t>e	LAI���߄ڔ�H������E�g������g;�g׈dC(ۈ��`��o���
��0��� {,����v�Ŀ��+�~�.y�n�	z���B�$�Wa�r�_/��W� v�Y�=9�:X#}�'�g"�� ��$E`��3B����X�n��?D��X�/zꋓ�q��k��Bqm�7�'��������w�Ǫ�p�����N@n4S��z�=�0v�
Y�y%��ZE�(�_����~^�,�R䨾W�7P�ڧ�9yV_��5�ZN`��S�|��._;>G�>	�Ipʍ��\����q O����m��~IO0}��-���<s����^�G�+
Ӥ.��R�w���n��Ș]���O��W�ԥ�)D�C>Aq� ��uyV�x�5it_^��AW��3Y��w�q���k����녻��'���3I�K�P�l�'v眚����*BV��_/�[ے����3�䍇t�<hIa(�S<nN��В�m�_�ΉA�����T�pw~��V�?J<�SL��cꢾ��X��Ƿ�;��Sb����y>�{��2�>7��I���f�}�.tf�yߦt�9��D�������ƪ�G��1��i��q�;>q���FT�B�C�z�׋9�/H5�Fw�f��I���r��%�{ۿ���]��3��� ��)З5���ͻ����|S�D~�F*��!"�������'�}�~Į�����d\!�)�Z~͝j~%=�76�Dd�^�����S�O#����������O�Z�fH�oP�B~B`��c��c�s>�~<�Lm Hzw<`��L$��b�m �#����pDzrږ�wZ׊��ߵ'��w��<�p����{0�*RAuh|t0T����C�[�����W����%C^z�6��"v̷ð"���q���o�~�ֶ���p��"� ��<����ɾMO�/x��a�N�D�����w��+���)~�ߘ����@���6]o|��3�̾A�!����|��dݚ�:�^̯��M����3/�<��a�:��u�߉-�����Ɓ�4/G�����~''K�gfK���O�g2��%��b[i�n��x�C���R�E4����sCr��y�9���S������䯙]tk��"��|�/��|��P����g�B���ހ�_O���*3���cw`�J�q��s�������.��T���v/(�O�{���/-%}LzH�v>��{!���7��1(�n�뀘Pg�1Vh_�]0%'�/�����.%����R�宯?��G���k�����Y�v���Ty��t�	��?�������GW�����s�*/hI���nm�>��!
�Ɍ͘���r<�j�]g�/j��iE.�X����<i
e�S�(���^��ٜ�͈&�����b�S�Q)f[���(�jL=�<b
//�;�r�1XW����~��=X�K��
�F+EL��$�̸JkzD$+�Ox�,�j�<E}9hJaXs#�`4��b@kgФ��X?Ic�^^_���>Fveu�~��+`r��w�]�1�匒i����`���d��&���ђ���P��큘&�i
�k~��m4�˨��M5k��\�Vy����ìQ?�oL
�@��[b�5�њ�S9JK��g��ٶS�DC䭃`��m�� �V �JXr+�	i��r�5��\k����|��sE��L<���~�dR�^�Z�d�2c6�$c#��!�UmX����˛pH~�NV���\�.�aeY.�hO�J�L}`O�a3�2VM3!͜�����G��l�0�Mj6s��Y��ݦ�M_��m���VwG�dT�f��i�#�%�@a1fl���%o�+n3n_���M�GƎwKW��MiQ�DM�v3��w�t	�����*�O 4��d�Yo5�a�ի,�[^�>vRs^�p!&�8�bq�z���FZ/�v`�;#��R��BJ�D�G���[���.��9���n���̛`�9��kgі�B�M[me:K��f4-�5��!(����s�o��{���	\�m���48�Nn�!!`ǀ;h�`qĦoHO]���X�R�W�A��#=Ya�K3�msn��a����IuDE��v�b{nчZ��2:h�ߒ9���N8�ա��zZ�d��͸�=�#ac�J�)1g:���0���n,���>c�D�um�{�-��\kS`
�R������qfT5l��?�>������>b:���G�ܥ=�`�(�6�ԳH��m��[����OM/�2�t}��
:��F��Q_$��Ɔ.at8�l
tpW��l-�nx
�$HN�eO�G�2�Vq)��4�M�<J+с�0�`�t}�pH��m�,׾�#�9�1Sb/*���ͯ �O+'ڦߩ$b�ŕ�z� �4�Q�*����,�\�1��/��g3@�a�G�mF:����䢠�<Ui?�[O�
=��Q6������}�pKLRQ�A�0�um�MǯfݖF�'ׂ���A�"��&��Ƥ�{"oJ̲܌�ms8�3���$�Q\v����6�;Ū֭�Y'��Oz�l��5�ƱʶJ�V�E�L6�,9"��C��M6�����|)`�V�%����ğ#�v���r�3\Y|Uj���9w��ՖxNI�v�G*��(4����Oog%6 �y6�v|��#��$����	F<x���6�'�Qu-�N�I�_��z�r�M'T�Y�n�:Ps9���l9o�����5�̌���ڸ�[��R��]D�L���j@P:�y����COW�٬Y�|M{Pђ��B!��Z+�/���|o�f��*R����x6�4��� ���{�F���7b�~]u�$ܢ$=M�z'���c�f��kri�8@�rs�څpE�M(�ٵL�)]�n�%�s#�ƩXLҪ�q�Y)��̔�Sy��'�0�.	
d��9�)3�̠|�iq�J�'iP�t�|���
�G�EV�lm�*m��^�s������۬�P�b�Y;7]��l��vy{�.QV� �"����bh5i+�����<R�l���`��
ۑ��v�S�t���v��L�Eȱ�Z���VG���!��Fvl�,��tB���њ3!Au�
 �tD|?���j��_��(_��5���?\wbl�S*�Ŵ��.ag,4?N����M��z '����<�
��e���.z~;%�����iuI杵�ve�*������ɻ��.��Z�1�}H�-=��I��	&VO��*�v��@�oO0儭�Iޙ�xĸ�h21/��������D�`���y����e�Y�Mכ�8ay�ݵ�35���ږ�kj�fʀK�w�!��U�=y\�ƴb�Q�;���eY�u���6������^�jΥ���#��椪��6R:.s�*XY*�:!�i�"5�[����40J��5����6h�aD�KY`�����,�
)���l�������^Y6G�b��F��s}q�����:"F���LԴ3������S����ŴW�1���ŧF��=�����x����[\���9�����ܦ0c�A�����-�[^~$��xE*��7$p��ӉuW���շ��\���7X��YZ���(8�U����ڨ�cC?taN�e=G�*� ��f��$�U���tÛ�����9��hs�{hK����%.��;�C���D���9��gY�\�-z��,�L��^t_9v°�z@K���ʙe�"��|���xOo�0�ar ,�����tZ+l�l�,�vS�sK3͞�Jn ��H�"�"��p9��,(�*|��yu��v�|V>ݬ�g��2��ᨰ׆���������_�^��Q��s�S��K8w��+�?�&Kd[��D)�t�F���j����
^<����C�]<��'�T����6���~i�Is��Ĵ����gC�>��RO���m�Z�b�u�`ۯ�*
�-�t}�<Q(��p�d�2����̪ܩ��?�SM�b����S�c-``(ALf��l/U\�,bC�r�
$�e)��;��X���QJgsI:�gc�B�ۺ�πyJV�C�$mf���˸��4���BL�Zc��m�=6'��?��)��D+RM�%�o0m2��"	��PQ�U�U�Ԫ�p'����bs�8�o�,�c�&�5�`F:����+��HW��۪�,���<�DS��/�cxP����In�Ƽ���ė������	ʡ6�S�Q�h�as��e����@k��\��
1+)H�+����^jU��Tz�k8�iG���"=zQ�S�%4U��~ ��E���*�܋i4+���	a+wZ�7Z_^J��ݏͨ�.a���U���8�t��ntb����3RpC�~)��bmI��h5J��hT*cS�|ZcLj���WZ���c]�tP*m��Ve\i���M�0V�ү�`g�RR��ie�T�!�XZӀ4��(r���f�-��~��C��k�+�Y��~W���ZU��ļ�4J�3}��� 7,V�:���e����uɊQ/Y�B����}z�	���I"��t��#�'�	��Yn`{h�`���Ӗ�k#�O��[N`Ly�����N��+�E��K3Wd��R��5f�k.מ�t�B1c�Qk��r�M�s�:�}=;�5���:�J�g-:���3��M��ZW�M9�J���c������ e��Ó|��0�P�u(Rr����8aOXk��վ���j�����mH-�)������������"�ݦ;��\���߱q(tQ��^��������O4;�ۘ�4�R��̶[�[�8n����#xS��o��0رڟ�����EdL��5��51yE%���h@�hH[�W>�����(��b��No_�@l3�-�Z#�S���ҟz�
�J����(W����x']���zb�y��7D�b�+�2E6���Raa�Gin���^�Sө�kϳ;B�n4$��c����;��
���o��}�I�/VP;ö�ˀ˕���D)S!��|���Y�6�Y�i�Q���iѡR�>�uR��3ȶ��]EkҶ��"�io�y��&(l�JE��v����e�L�V�**g/^�������o��K��׻CVD>je�c��ж�(Ԣ6Y`�+-��Ryi���C��gj�[GL�\))z������k;f����6?���fYv:Գ7��v&ׇX]!�R�E�ʶ6ш��J �|k��<�h�Y��$�o�y��Et;/��d?Ԛ�N��`��Zw���j��Q&8��S�_dw�,���*����A`}���Ls���z�@S!W)y|u[�!n���rf�E@:�B�FG�~�CG�@�ƻg-	��7A�i�=.i*V.�8�L(�Xh���;���êp%���G;)]�]
�q�5iC�<@�`���5��I9�g��b=&$ �l�<ysHō�L�9O�8+�p�*���0�kj<p�osU*��И	��rT��	�[�p��*dQ�(sәp��h?����gVC���o�W�s�ϙ�wG �b��u*D��$��H���W\J�f�JϜ��X�h������#h��V��.*��~Te��[���O����.��zUg;I��h�	 s��u��+���Kk�:)���1Ft_OO��xMI����p�Ũ���D[���r	�S_#�Дa�˟�+�ݣ^�	!�i}�$���ΧV%���N٧pC[i(�<ֳnVե����'s��6B's���ÖB
��kX�OR�7��P#Psl�_y�P�T2QP�:I���U��u�M&DKJQ�i=�D�b(�pw�!��K~n��
�E�Ø��0�=�[��,-�:��xS��uZ2�5Y"�e"� �j��MGF�Xtf`�� 0��!D��@�kV42-]�w����P���6�U��fW,{c�-�F�g�HLVhR��L� #�LJ�Ǹ8!����R�<��L%7�K�zcd���D��V�Z�'2��Y��6ɑ����ؤ�|q��D��g?�(�Ķe�J*��\�p���,�5i*���
}1�������QڗɄ�X9�4�,Εr��	:[hTH�$�ۖ|Fq�')�=�Է� �'���:/�Hu��{�'��?dC�<����}����l�'��l�f��`��vhu�{��(ԩ1�wಶR���¿�¢�#�qv�N�Ӧ)�H��vUv6�e7��k鎄�c�f����ì)ttt�\P�BQ�D�Ȇ�݀F�|Ij>������T��ԥ�o�HE�i]y;=��D3�v30�G�k������z(��˝g%
����`g�QsQ�'5{0��:��"ժ2��T+(� vz�ڕ����u��"`��)�so%��U8����H�x�r�z!��";?("/��:i?��W�_���G�ͥ�Ʀ{�=fuL[�T���-��@=Ug��݌�@��1�S�$V�꽋���X�#���p��
�;bF��硒����_ۦVLCl@'�2�b���F�Xob����|_W[5L=���b�|R���B��U���\K��5V��,�Jo0����2��Wt(�zs�8�����+�m�H��c�rA @�sb�݋�J[m��[0��8c�`x�дf�
s�\>�ћ@)mO��m(�Ц�O�I��ͥ���T�ޘSt�,q$r�����U��]ѹ����[t�=툫I@�����D���+��a%�E1X���p|�h�	9�f��
9�ԩ߸�\_z���,�eU�v�F�h��fN+�.����a.}$QQ�+q�I�Z/m��!�ɹV�]{|��c�+���N����R�1�*��O�;�F��)t������_5g�< �%�21hV��5O��*3"�5<�N�\�w��B&��{�E�=�g��^)8[���CʦquF{�Mw~.A�� �d1������9�+��C��~���L��AD=�X�*	G���0���v��<BzA� ��z��ڡ�[�wc�3ULȭV��=�CcY��A�s�׀�2���Ҕ䄠I���U0�HO�_nu;T[��W��i;{��4����V��#p���a?H���'X�Q�����&Ū���,T'����%TE˲���_h�� ��|��&��l>�?Y��d'�����C��$cz[��!����Bʯ(���F��Y
��;��7�&`��]��m��ƨ��,A�,�l�}hа�*�ğ7o@��D��ee�K����٭�-�Eއ�����D��k������Lǖ��/��8�r�vee�|I7Z�yC�ܝ��ҡ3s������#��CΕ�yD��<S�,)M�ߐ_l���D�Z*ʒ�	��Pc~'ޔ�em%�\���]i����!�������M�Z܄�~�_� �fH-��@�q��V�J���´,�����k$���8.��m���Uc;/Iܘ��^�^<%���(��sTP[;"�J��?�A��V���J�<�d���i�
 ��b�6����Y��&3�U��	��7R����-:'�V��p-�w���m�yw�VV��PJ_�~Հ.���yJЖY0b���lu�VU8�?�q���a܀H����Qݨ^L�=�3��p���J��Rvs܁��(7��
��k67�&#*S���lS-�4�J�ְ�e&Z�"��ҨLe�ZC��U�0�b�˶��T��<�F�f�v T͍���W71v��ԉ��$�jb�"L\��j�����'-�-�]��UFIrBO��-�����gC �N��������r����fF�n0|<�|��.;������G�Φ���fZ�Kk��u�1z�S�Y�ERG�g���˨��jZ�BF���F���9Z�|�����@őb*�V՘zj&�ک���gm:�ː"f];U�ck����z�IX��1� J����ΗB�Z�&d��
PG�s[�Z18$*����eU,���*���IѴnB^#��M�H�n����;z��nc��c����K�5��}�t��V�Q��R{ה��&xd[m� y#`ԣ�-��K)�Eq��z;��`�	X8�~����6��:bz�������Ҥi�3r�\x��@�T���T	0�H���=B[�'��jv��\�٘I��|�A8�������%���@��Z��[�ꌝa��
#ߏ���f��<Л �4�#���v&���r�WC��}	�f��G��y��N�DZ,_��j�v�Ԅ��J��<�^�?G���Ij5����%��������Рg�Pj̷�&g{���9�Ģoi6�s���0!���֏B��]����ƿ��և���~��t"b�Y��V&^�z��,�
t����`{y�Cg{�)�䈩m_
�}J�9V*�(Ğbr��8@��{o��o_�7:�o7�5"GR1Ic�>r��&��I�&����.���3a��k�{��,>�{O��q}KԵ|v����w����2.hժ�-!-�$�O�(���WZl]��pN\�^�^� (pC|WYi����'N�M�����Du�s+2Ey
���JF,6������cդ�]��p,K��W��]���fA���wh�%ɹ��K��O������]4�}7&�{<߃1��1H���o�w���0�,��/���"�ǯ��X]A���������O��Q�ͣ�ک�*%ص�$6�}�{�|�g�`+֙�xD�l^>㭪RO$'}3VV���!6�兩�8t�*���o�w�����?ѣcC���gO
�>���W	�QK��5�~��w�]� "���VA���<ۙ|�����Tmn7{��o���?O�}�7���m��h�.`��?���G��敼�	�茜7}��3��.�5�?�6B��!��Q� o���?6�96+�)��q�9��Ÿ���b��ᗿ��G��~���Zhd��1T�n�"z�w�sI��'���r�k���g�֫|�
�BQ��5X.�K鈦��a.R������\^��_�x'�
�V��c�uY�:7���ElB�N���c+�~��C`O�@Oѐ�/��D{�k�ҡ��
!C�=`"!>�1�R����Ǩ�1��M�#3���+�D)0*D���f�]���*'a�T�����eb��?��j���þ��ޓ�~/�e�6�% A9(�&�H߭čl��? T�����{�)�8�e'�ϗas�@qz�1�?�u��i�$��UV����`nm��t��\�熈ЗBe}�ql:?�D(�2���4	�[}�3�~N��uX��K�ڦ�p��k��?P��n�ZY�k4n��2�D��i:��|7KXqb��5�|hl�0��}�\n埵�X�?7~��֖GM��RJ�ٓ��Ζ&<��8��ը<�-Vr�q$����[�+�t��d@�Fe| V��F��7ߎ]�JH 
��'�N���|~p�ʼ����dR��>]�rn�����l]�%j��ӟy�� �.�!k	��Y�֡�?*wu�8]5�($T��x��j�%Swl!U ��)�+*1y[1���y%mr!�)�dvZveh����c_mS<q���6��x�iQ����}�1��R6eH�-.d9Q	(o�,���xa헆�P���a9��fu�jƨP���֖i%ڨ_�}�'�\�Q��1/Uoh1�|��8M1烙Sr�O���;WN{'o�J��-Qoa�\4�:��U+��Z�ӜZ
ڠ��U:h֑&�cI���i*m��ᄊ9G�B%���3a��ҕm�JRg.%T��rQ���s�_���5El�eo��Y�4st�\�E6b%�ZH�M)Q=]�1y{t�� !�/���Sa��QY�57���t��m�TU'�h�t
Y��ՙ~�(Zev�t!�8��)���l9[���`~���X�;n��lN(F?@��ښ�Tpg��4A.�����S��3F%J��m�u��04�������ji�Wm�'��)��,��L��f�����t�z��a4a��y[��٘�\��H��cj��e�JN���ۏ�_�c���^E�͔�S����	m��b�=F��;�@��`��rS�E<b.-͊��e��i~LJ���q�v�J'XP/�㦢�����Q}��bB��*+���mX"�kh�<� ���2U�1��o�{����9�`_�87�,)¹n���k��F��3W�z��c�u� KLNһ��R9t�N<C�;�E��;�R�R��YI�U��m��}g���c�۳�w�^��Zm~
��������I����aI��⤕=��	�f��9N[8m�V_:��֒M�籨��U�(��<ς6M-g�J���ť�:��w���ԩ��U]:��#I+����|*X'�7p���Ɣ	�s
m6W��X�nT��DX1������*`��ܘ�§E���)8d�UQ1K4yTuM������Z͋0'{:ݨZN��� ��C�n��<5�	<?��Q�U3�'���vub�F������u��˙��Jj3zw`��KR6Ӹ!Ggs�&�f4f�%( "��f9H����� j��-����i��ug�j%�"�����g�֐�=�nx�(���=�Dy?%V%�K"��C���fM�.�o!�U<�Hi���Y-(���I/
Y�����4�l�еQ�-eb�i��x09��H�0�c�VR���,�9.�B+0j��xgλ�6m��95L��]M�bW�����
^����jnt�)<�Y)裧F�)�4!W&�2B�uwT�٩�ɽ���T>l�<�]���o�[��� �&<�VE'� ����LMiIS��	���C���[�&�N�k� &^�wk�5 u�ֿO��C�fQ�.���t��"�M�N�Wp�LT���=�l��9��!�U���Y�SCǱ�	�D�+3�9��IJ�1i���%N��Yͺ���r����6�旑��k�-o����3߼Ò�nSX�dM�3"�Q]��Q�'4��I����&��H�y-p�5���[�+ 5�%�j�xH��&	B��Ң��-����X?_���ɷ�j�S�˫�jI�pv�.+��y�Z̞C�\)w����c��=+;E�H((U�u麚MJ��<�b8:��Y�MK<ݸf��Ь�X��|�ҘEq
�J'㒔�[�H퉂Hc!��Sf���˚�Q;�e�cBn�\�p6��z��p&8�ì4u3	�!NN���8�hʑ��;1qB�$��ɸ�j�D���e� <S�U��V�j��UД6�n�R���hզ�E�i���Vp���7 �%kI��g0�{�\]�%�#^)��(�:�ͫ���*�X��G>�}�豼�t���}�ᜲ_�欘H
�v�1�*��I+J�ٜ�ɤ�����O3�j�s��D�V�oN���;l�]9�B�N`��t[4=�M;���6����]����*�/̣p��|��y�A�W&�1$�p>o��2O���1}�y�O�>��s�_�Qت�s�Fz�D��6hG5>k�1�s��M��~h���� �y�
�eu=3���Ge���T�w�{<�Qo^�W ��A�L�#^�0���Y� ��4      = �{Kq���Eq�/.�{���RQP�����B�%�R/.�{�:@Lf�H   ��+$��)�	��::�`i��_�X6so۴�ι�����g��s������b��9�q'��r�Ŝ���{
/�l��~"�1��   hF ��n��Y��ֵ����$>� ��@��BQ@��8��I������� &�Qp!�9�f�΄��-��5��&�3�,���e����m��l����v�K'mM�,� H�����%�t����t��	���Y���k��W[./^wq?�}�N��m�-K�k=�̈��g/���ewmm���������d�-]����g�k���=-���{��8��ۿ������iˬ����[|���%���9�u��g�_/+'(����|>��͎j]��2��,c�-z��g�f�>[�hQ�#�ތ{��پ��Wd�����u�,w�L��;;��"G��v���}�_\6��_qw�*p3��{501���@n�"o��6���\�����E�m��d�n��Pt�FA.��`5�?�6'�o�W嫺"ތ���R���n�����G���o��~��$��}�̈́���>��l����_�Uؖ��x�?�	�	�ư'��s�?��z���~���'���_�Z���RE��!� ���� ��q�9�xl7���R�<��(V�HC���֦�ذ>(� �����c& *
�$&*wc"������$w��B��?j��v>&����!���*��xQH���.��<-��jq��'?�:ܣ��Mfr���b�wj{��U2L�6���q{��b]0��s�7���%)�Ī�i��%31q�Q��r����%�{:cC��8�$ݹ��� ��j�s�td�}��q/^�D���v�� �+n�וZ%! �t� �N/ � ���i����щ�:0ߟ]a@ShM�3�չ��fb)�������v-薍! x�^?����t�!�/v�%vX9!�w�^�Y�@D��jA��͈펄u��OqevWv�a{f����q��8{��|��:~��^��]!	ݞ;�?�U����i3��0F#���!��2������jȵ}�D(;J������-��mx��	��E7��"-$�}�A�
� t���A7�b�����m�N��T������MjweM6� L��p��S:�b��0�#�L8h̗7x�1�v���+G�'��%�(k9�+%@=N0KlC����p�I�������<+�7J����b��=o�����������s���������L�C�N�Z̧�}&uK6�
T4���ohyS~���s�Q�)�S���/��"r7L^-͸��	*��q�4�=�Be8	v�>�K//"0�;�je�S��-�.w1�-�n�xCuxQ�8��Q�Sv�b:�>7Z*P �D7����!�U�QP�Ī�%/�l��p�k�u$	���g�����q��\�wd�8��:/FmE���q� ��&jS9����5���nH�b��䒋��rOS5�����v�%�^O��Z]�Iʺ����qVP�5�7�rM�γ�(So������eBQ�b\T��؝L�����8'�M\��ŀ �3b�K]��q�q1��/Sځ�>H�Q,�f)(d�bSP����=����p]d�6��3�D�<P`̛�#���a���=�9B@�9hDT���A[4�}����(��"���:�c
u�p�
��tF�Q=gT.�(J�J�0�3�	M.��;P��L��T�".C#�c�Q�3jg�z�������,찈��D���.���c� L��rF��F��_r⧼<�R>��i8�n�5Pt���z!�!搻�YU訦1EÄ1�[ʐڜ'�h���ܤW%,(8�1��{��=,��1��6����7���o)M��ݾg"��7a���7wd�4e]������D��yϼTf�=+����eT����s������T'7J�(��x]�ď�n��;O��E��f�	܏�$b]�
���l����ԉ��2��`C�Rz�1]�xpz|SZ�"�W3��O7�D¬�-޽���( 0^$Z�&Ș�Hͫ0��sV5��Qm	M��)0�)���М}ƚ|ҥ#/]u���c��`7��{s}��?���+3MD~R~ �����	8�k�5B�f��um�t�:���qxN��O�9�̎+�Ӹ�)w��bW2$<9H��'�BL��{	MMFi�w�^8x0�\,��#�x����p��g�t�3�P��%�g�Y*<k2Ӡ����s#sD�Q�y�j5��-��	�5���y 7:���Ɍ9u����n^X��99��H Iu/�K�.�K�p-��ԃ饈�p���e�0�&wA�`�K�/��sV�^���)p �MD�۷KAX����������:��(\���gJ^�;�vd��j��.		�zQ\Q�;��Uϧ��	n�{�*,2�lW���B��Epm�����sy��X`#S�Q.��ҊݣN�aKK��Fc{7����I�U�q6&U2����A.��	7�r�ݵ��M���Ma?��4�r5�bHk�+:=ɭ�h��N�{�B �m�:G���WZ�P�����ǶY��#1��%M�j���jNU�❍�^�d=|a�dm���#��J������P�X�#�� �V	��U@��o��$f����Ѽ�p��A��K�N"y��֨�cJh�����!�ߒ��p�j��\�<A=�a���'}	��_:r�%n Dp�M>JQ@t�I��I���ˈ�ƴ�'~�~�	!5i��y�$���V�~���	�>��N�������<O�����.69m>#�˱4�5t���ߓ5��k�7f��ޥ��*6㨝ð�A�g�-5��kg�3�M�e�g������m�9����1���`�{d��z��Fx�oпX_�d2 c:���������������C��V����ɼ��;Y�
��u?Vޝ"���Pއ���h�z�U|�W��̙��_�}Z[&��^y����\���Ӽ@��eB���5�^�oRi�,kM�~��k՚Oo�z/c���
ѥ{������4���g~&>�@r��<�tk~�|���-�!�q�e��f}��t����`�����K�K�	>����	׍i��wk�@l�]l@�ϕ���z�ʗ���R2�w�j�d$�wNq��S��o�;����_�D����Y0�a8������y�3H��R~�`]%[�m�����v�[��s!J�!E?L�89?>E����{�z�������z�3ވO�����^��l�o��=����iR��(W۫�>0-�a��y�������߃�l��������@�W
x�(����Vt�����gu����'����(���'�e.6�~���i�q��O �l��=��a�����2�S��_ۋ<���xv�˙��r�}į�n��U�_y�L���b���$�b��?�)�	Ε���/������jpz׿��?�������}m�ϋ��g��+8ʟ�:�6���������{����hߤm���$�V��������k@c��//_�?�����_�h妐�?�?v}��"��~�l�D�}�W�|f�?6�Ed��Q~Eʋ�� /L󖆙�1�2��k��Vx��7��ݝ7������s�x�G���>E��-���2����}ـ��� ��.l��W-~���`��So�7�������e�}�e'ӕ��w�^�?�_�bjgn;����[X��/��g�F��U�vbGv���S�o���09�`x�nm:O0�>m�0?ty��>/�!�/��ǳF1�6�j����~���u�2������
�\������I��n�w!� �g�Z�Ͻ�Ф��+D�?�����J�@|g��e�߳�=���������~�}}t��5�>zߖ8��������g���d?�=�8��S>g>���'���~���X�vvf64�}"��~�Z��q|��K�p�;a��)�2�'�O�z����_�Lv^�_��T�1�m���j�'zz�|��/�4�zA_���a�}�A���C�7���&��q��zCI[�F�?he����> >B��g�N�E��_��]��OW�<Sǈ�2�����]�I�P�?E�$k����=�(@;�?^U~*�7l�����+����da��/1�|����#�ol_�����K��>�'���~���A�]Oퟓ^H�~�+_���_�i�J���Y��`����A�y6|�������
��8�n/�nxP�^?-��L�_J}tz�ڞm}��������3\��}y������9�O��ߠ�Ժ�(�?�����n�RO�o�*|dc1��z��f�?f�45��yK�\]d���m�F�����x'��|����V"�M��?+_����eF�ϻ���~����I�}���l���aӗ�e#���=�;�< ߾���'�*О~ϐ��2�6}E���!����I��X�������˔��N?�{W������w�S���$�������}�r$�{��?�6��g�?�g����B��;�^�Yh�5?�w��O�����2��~p6r^T��.�iz�=%��]�1��}����oq����op0�H�?�����+�fS��'Y;0����������_Ф�}��{��O��?������o�V�����c���o���-��;G?;��6������=���_�u�`�kW�G�ÿ�C�����w��}��~���On���_��!z��Ix�?^�������k��s�	>���?���H�S |������G�vfo�XI��ɸ��$���2"*��l�B\_Ҭ��Ϙ����k�>�7����_|&��W��l������l,�~>�'��}�~&���1�u��VSP9�́`?���\U�����B�����o& 鲞������L������������N,=�B'�W�*�tz�]�����J�\�s�C��k�����������}�F���b����j���c�Ol��d]�z��a?p��4�~V��HP��~�~��&��Ux�e���y�����?믏�k�w��?�Y�+�����.}G=��E��h�_i=�zH��0Q(f[!�{�.�*xS?�$�����GE�v�~�\�����w��9�
�a�}t�T�z}�N��ҹ`�C�o�ה��+�e����M�������_)�ge��O������-���O����?ο�R����>�_/�4��������~�q�\ߞ<q�K��� �a-
jHA�/��]�~�?��������͋���
RHA�/�Z�Ђ�������/��^@�t�����;�}��#�{%������O0&�f�s��SWL����{�v�c�dW�������WM�VY�p���;�|_o�^|�9I�>��?̀a�W�����%�>�����/���U`T�A���þ�ݷ�N��o<�v �do�E���{�3�M���ɣ����;k�"ܫN }�B�T/f������?�}�~�_��x���"���3h����z�^�B�/������C�q����t��f�,hV���r�m�X�j��:)��o$�i���R��r�Im����fv�� ʊm�z�H/{���we�\��ax�m�\�w++-ŎXU�-:�y[��EV�7^��H��	'ε9�4C*N�T���Q,qh痹B����R�D���9�Jg��>��O��i�Z��o�\���Mҭ0���|U~�P�2�c��	8E`�}�j�t�%ެ�8�Dw��֊9x(���p%_a�(��@2�^nk��	/�BA���m1������0LoE)�\���46��A��5؈��v��&v� ��4P�
�;s�XlE�qk��V*r�F������4��N��h������fΊ�7�:���}�c|ʳsh����p�l-�V������UV���0�,��Ҧs���F �*�H�EAk�	rX�+����#n�r�T�m�U4���c�9~c��#e�`��0��`�c�O�x���S0j	�������m�k�lin�L-��aW7W��QO���t%p!6�p���׋��&vg�o]���Z�:��Q��[#hK3m��@�D^Jd襯�JQE�I��M�&ô��uGz��M���#ŕ��[�����6�IE9�#SaՑ
��S�g<#ڄ�=�G�>_�T�B`������¡	�m���f����	��r)'1�ԫ<[�m��[� �3R�<e����Qk��c�b��W��M�'O�r�;�lNM����w���ŵ���c��~G��57V�H8��X��NII��f�[�9�YM\�x��W��͊�H�F��U�r
p�]���FJ����0[���\�ru���詳v�]�������7�E����K��GY�2,hK�!��"�x䮍�(�:e1��[�1՞i�N��\(��n��Q/$��M]b�"������p�-�m$!iHl�5��z5��4Ƥ�NIBh��t�(����JFP�&#���4�T�8rM�)�̶h3T��	o1�r9N��^ś�o�?��x�N���އ��?)��Rk�ôo�7�@�G�U^o�`#CM�ʲ��� _�vP��S:����}U*N���{����aQS�E1@�e0�Y񂦸���*�mRІ���>�q���:]�i1����΃
Z�o��
8�N�	�	����"�j�<�`0'`i���֥�y��n��eB��x��&�Sڼ ��&�����v�q.i��xHæ<:�-N~����x+��"zye=���D6�3|��¯��5g���E ָ
Գx����[��rohݕR����Pe�#4敖c9J�������4�I�qJN�+/-�&�y`}����k)E�$(Q��[�7��ڹ��"�~��~�s��O�\"nU��Z �6��c\��7ߖ��C)X��j�װ�SI����U9�fpM�	�H���;
�2�8��@>3�.�����K�(�u�>'h���޴��6\96��*q��y�]�)�Ε�s�T�a��ܼW0(���6u}	0�A��+b����]p�M�n�R^"�f�Ss��kiM�����s�1V�KӀ�<�yZp˯�-�ec��ݹ�[By]�]	�d��v7��t��|
����~��l	�PQ�9�����mK	�d����a���xk�W�3�<ۚٸ:Z�s���q��D�fPxg��ѣq�P��c܀�����\--���qSt�|	�3���K�d1�$�N�����s�k7��-W�����s�@�l�R�ow�<�d��ݨ��=�q����-iZ���Jb�֪��2At\����/ϸ���J-��I���S��Q�r�lYt�XmsOA�NE�\*縶 `�<Ã��������:Tz���y��di�b5A�Ⱞ7V`�'x+�!Ԣ�~ݖk
��Bϭ��R_̶"	�g6�\y��s�B�"jd�W�U2�p��]!�mSb����.�U���x��qYc�Suر|�NL�k�����᷶�Y�I�:oW$w��ݫ��v���b�_�����n�7Ѫ�oͲ�1�}`e/;ͽ��SS�Q����R1����1 �� �=x�|�6�W�ܣ�x0	A�4����-��f�޶�7Jd�$8���Ԋ�q�y<�o~?~-/�K5,F��?Њ���С�^5%nTwPy�r�=���oc��c�����)�]Bh�nh���!��t�#NOټN�`�l%��=9K]��Q2�M^�mP\�	%�.+L�lY�θrT*��p4��$4:dLUg���9���������]�X6|NPZ���Hq�Բ��f�g��\n��	2z�$�N��y���L�@ļx`f����,.ǳ�5�t��GKl�i��7[ic���%v(�8�;;����ήwᡁэ�Fdǁ�ydY�}ܵ�R�'ns�.L����K>xx��i)��/j���7��m�	p��^xi(�&i�W�Q�{ y����X_��z��`�R�4/��r��q0���[-�t���6�S//��\���1B\�(��ne�B2�AqF��.C&iS�6��q�1ƀ�@?#r<����'�v��Fx�_�&R�wE�(���PD��6!e�=b$�J��ːN�;f���тc�Zm�B�0N��(�ھ���UKX]�Ů���d�A�|�~�&���4DÁ`aE?2d4`A��s@,�2kl&A2�N�<�V�鲘�Z���:iZ����־�\��|`��`/��q� �����=���G���U64~N�\a��EFK0�6��ХTr�<�����P/��A��JV����m#a
��00-�7M"K��MJk���*��/p׹UH��e���w<�Q�D�%�Gt%̢06x�yM����Y+�#��5<?�)�:ѓ�e� ���B_�΋�e�����&�xi�VO���	�4�k����&������9�w��"KK|�ng3��L��N::�#���6�4��LͮC�j@K�13�-��	9km�9	d���;HDE8{����0�Z�5B8I�̶(���u-sZ��Z"�K��ېVB�������i(L�i��ˀ�
"(e���5.���w�""8�0�"�+����?J�Ak���+��r�Y�X�#� $�Y,�J�,H��4y��"G�(0N�]4aԱ��#���	�Y�vĘ�0x Dk�jhܘZ�՘�f̣��dЕ�#�7��Q�u��Ǳ�e��)��f6�ɐ1���QQR]�}<��6�= ��UD3��F~���ABJJ��D+�%Yd ��a��~ū0�Y�cn��gQ"5��,��씢�k� ��Y+tR!g�6�i��ːr��2&mXE.�F
c��.f���a1d�}v.�N�dE>F)'ղ^��71��9�	�0��Ql5�w�\R)	����5n��I-��߉�7�:�e�p&g�� 15�]n�� @[��%>�X��^�G>xX��N>�G����L��@�J
���R$m��U����%��j=���K��o"�G6O+�½�i�^t�gS�s�v	�Y��'��k�=\59��5��o�hu�3�sP�	�H�wjH�DI�%ET֘Y<	n���D!\�_}*�=ke��$�[e�2�n�(>��`Q��_�Nyg1h�K��
@�3{�DF/sG�K�n$l��	6N������7l��Z̴vlH���u?�6H�[�T{�b.�)�J��)"-�?K�ȏ��OQ^�����=%
���j�E��`�����*��-�~�1�_rsHa�K+F�(�́�wǞ7�
H�[��P)-I�MT��g(u�c%��N�L�B��|��w�I��/e!j��tR���	�ҙz�{Ŭ=YFv��+A�̼D�ꎃҌʎ�xb/J��bm/�
#q������&��9��N2�Ft��dT�?o;,$�E_23$������PԤFapj�g�vO���MR"-w�x.V�%�
U�SRXk�P�����4�����#Z�cj��9����.=G�Eөt�����9�h ��_�o
�Ťҹ����
��
Jʯ�o�j6�6 R��Ww����N{���,p݅Nn��+��n�벲�8����N�1)S3��.��tf c�eԁߕ�T7f|��m4ƻy�|��N,�e�ss|�'�[���0��M�u��h�]��MN��"���w��d�Ac�8X<\��Yu��&��>'F= �	�*�g�C�ܵK#Zr���}��i��\�ny�0aW{�O,>���-�֗��՚���ϟ�H�����gThg*����~4�
F�j�QV+�-#/�����C��3UG��=���$?���j{y	�s!6C��T�FՌ�Q��] ��o�n�'��sn�z��4$�����7[�rs��ā�a�zH���L�V�V$�q����4�#�E��yCnj~g�XK��ƍ�c�jk��N�7D8Gƺ��X�������箃l9P��)5�}v%B�w$��q��ed�U�\��h��CW�l�ӊ\�x�g��2��;F�=�7�MdeO��8m`4�/�K����hTNf!������� w�Tv��#��ͩB?�u�n���\)G�jo+��" �dUq�?��kC���Ƴ�Uwp}���v��i�h,f�̬�H܋+H��
$���ez�S�K�Py�O�} �!�-��g6|+�����q͟$[Ya�t-�;Gkl�ԫ���K�������j{,fr�AGAA�6��e�^�ku�������j��E3!���)��j8��A��/`J�s�Hb3�|:B���0#W�� �G�]�p7�n.�ɭ�-��+G)��p0�'͵m�6�q�����$vy���M��g>���rVYF��:����U�����v��VT��WO�L��&�=��\���+�wzz�ٝ;�j���u_-�v!�ཬ��v�BX�9����lY�n��6�$�D��LO�/�YG��X�Խ����0�{�0[��Ȼ�ay����w�oe��|CU��Z��iu�ϤX��JHl;/r��L�����aՎr��"�kDxw*C��N�Ac�F�H�@Z%2L���.�Uu͏r�sy�a��/������`���0��r����r$i��l�j>�~x
�?.O9�a!M��w�������NX�� �ar�K�`��,v��V^hy�]gP��_�ї��.#s��Xbb�j���C+c7�B��W�O��X)�pj����C��p5�X=q)xn�6��kJ��AѤ���J�k3}�m7������ @/��:	��icՇ �Ʋ.�Oc1uj���MR�W�X[[�$s�gX9:Ac�������#�������C���P����$�uBh�_�^w�����=E�ꃨ��h�]BpW4���(t��q}�{�[��
,�~pѿ�՞!.��;�$�R�Ը�nUϷ:��#�K����F�\�D�M�-_��
�C�Q���*Q�3�<Hj����;K����s�Ũ��S����!��lE
~�;�X�=0xda�)�����A�V pE��e}� A��N&2~�q�o1���
���
��Y��g�aX{JY��!�����P8���/W��H�B�:���X_�y�ԉ.�`C�{9�9m��x@e-��q¶*$Ax>l���a�����iU ��:Q�(4����K�� |�yV������{��q0��X��[7ܘ�6|R��X+aɴh���t�V������ ,��D'+������spy��k����
�	��e(���q3W�����/�S��v^��vdJ�� 4wY�� p:��I������C'w�7P��ES�����L�90�?��U���0nc)J;��hНL���n(��g�=ِ�Ǡ��,T�����qD��]�9�J2g�iztt��[���8^p3�����88�1��-㤕�"�OLZ[@ֳ���`�R�O,�����1�	�W�D �ܶ���9�l��Ξ[@ 3I��b(�),��'\�k<<��CoI��i��J���bW'B�j\Lmk!�ɶ�|o�'ݧ�C��}[/Z͛�u쇤)�q��KT�$���v����������L�m�^��,v_
|�ȭ�`�����&h�ыI^s�'��k��r���=ȁ8�c��;y�a̍:-}(������u^l{oG�lP��v�ƫ�8Z����ѡ/#ٽ�?7���P�@�ХpM��[�h@�x�4���-|<xE煱Վ�X�#�z�z,����%؋��s���X��N�����%8"�34Gd��.���S��Cs)��}E_M_�+���ȹ[x��a)�bl�#����K�bPrg9�4���b�Wp%1�,�7!<�����j�!�A�y��H[n)��cB��J����n/ ���O�vk�&H\�1�ɮ)<��$�%�s�2���������v�`x|i��л�2�27a<�g傓q���	ouک�5s3e��;���LT	�xW��%���L�QMŬ5��X0��3Q��+�Z�;3���9�BF��!(��{P�X��=@R`�W$<.� �f�;@��Z�AD$C%`�!��iQӜ�����
A�_�)�TX"�O�h	�]͇v�X�4^(�*��)����b�Io�F&J�6q�K��;�o���ё�Z1;1���}�o�GGWo�jT� �݃���b$��R���Q(�R@�����o0=rY�jt�V���vt |sz��+�������_FFa\<D���oFt�b�'��B(�����r�Rv��$�p$�C�x��)3M���_X)�zU]��'��h0�� xh�������vD���R;���e���^���V�ƌST�H(u�7�*��!
�W�o:��q��@u�#Dz�}I��K���=|ȹ��{��¤T�܌�V[H��x�r�����e�-�C^y�lxc