,݁����3�h����.�2�)j�����J.@�3���mܭ��G�8��["G��^���WRa�G���w����e���~�youz��1���~4(����԰Z�[�:�99�F��KWe�k�+
�O�����x6��B�hAF�VY��BUb�9OC2�u&Y,7/1ԭo����Q�����������`�c4:�S�[
�F��W���X��ܯr;�梴DuO�H��@ml�IE ��!}�!�?�`_c��i?��=/^��dͤ�'9.�x;��`A�`x���:k������
�Er�w����J����C:�{���o_򕗔��G��͒ո�0�Sot�%!=�3�WP��%5� �NX��'ڠk�\U�����P���7Z��g����Dq�� ?l����zy�frU�W*��3��s>��h��[{!�����5q�i��㛇�kBi��ycke�צ�h+՜c9�������n���˔�w�F���!/f�
 �5���q�`�J������x��^fV�'�`�b�����UI�tT�_��-�
xU���Z�Pe�1&�9��l�!�%B
S�_F���]%̟3�\��xW_�B����{{S�G���(F�>"���aI��Ĳ���ޛ�q�t�_�B���eOߩ@�.�d7�U�q���I,�0�*�����H׷V	��B
���
	����x�gۏ�
b
)w���Vu����Z �x�l�Đ��d�y׆g���4�H������YV��W�U�����-D��;���m~}��w�Pȿ��D"Q������|l��+����|Ѡ:�_�9U��7�8�UI�3�J��Ɍ_�i�_#�=
C�~���"Z���Pl�~ 8�ȱ?r8�+�]� +�; ��l� 
�H%�A�����`�%�T6��������ӪK��*��ڹ��2�v���Ϣ����L�w�q/ow���n,P�d ���و�藊-�e�	
�ؤ+�H�/���S�ȕ����.;�7:2�S]�\�Q�%>��͂��ۖ卛��>h+ V�g,9�4�7Tu?�P$_3C����s� ܢ�����&�J���?�+�U�Nd�J��q������ػ�{p±���"����#��S?G�xu	�Z�Bkv��L�4'��͉�@p�+�� 	s���c�'�b,�P>�Fx����D9�|������rd�%_s�|�p��gӭUU�
�bh��e�*�S�ؒ:���8P�w/��^���{��>C�L9����5�;��m�������{oHm��R��#����m���$�����L��w%)�LM�l����P�c���_ڢ]'LE�њ�9��� |������6�5��-�����_��-n5��9�8e�O�&WO�N�݆f��&n�z�E�T��;?�`i܃�.�]�zg��pE�uA}���oO���:��a�s�`�aD�럓9�_8��y��v����j��e����	W��eb(�o.h�s^���;	˦�x��iϜo`���̭3n�&,�����:!�	h�1#�YV'�C�����-�IlV�g��l��I���)�9�}��Ɯ4qPk�]&�i��^�ܸx�8��i�����n��; c�N� �|1r�e}�ԦU�6��x���R��߉�����S��n;�B������/Ϳ.�~e	A�7�T�G�Tا�<����LrReU�o��ς"��#zw1Sq����o�P"��%������i%����K����
d�I���*��򦘴�]!U�r���E��C�V�&��S�WԨY��n�jm  �]@(��#9W\����5>�G��]�!T%u���vyx���j�6����y��i�[J��[����p[�}��7h�7����z.�B�B��7�P����M�G����m��*q���2���H�+��=H�b_ʅ�l�0 �Z&�C3�Z)���r_ h�`A���uE\��}�	9����^w�t�[U�;��o^�̚��x�~���B�ʟ+��G���}ط��Ex��u]��2^?E����%:�#������}�TR��Yה�5]'��tU�K)��Ħ�~����q��∐��wm!�wD6F��\�3yQ5kC�ݩ��F��6����J����� �����G��l�� �42J���K�<a��m�I���T�8(�8�ymfk��+�ǅ>/m$�V_^����,K��0VCOwRː&�7b�����ZZ�k�s-z�nQL;Gz>�9��;3R������2��=�G?b�\,*]���=:��+�RP���#�V��:)ۃ��̭	�;*6��T��u���;+>\�PX���V�z��nr-�t�͂�()Z�"�[d�Ԇ`ǵ;%� ��"���ef䧉������G�8��;$H�N�p�7j`�vU�+$b����Lm&�$�PЫ�7��?�Z�h��jz�>�e��~J?��iA�|̔,��H-���ӱ���[;N�@���;�ت��N�q�X�^��&6l2<>g�dޝ�m;��vՔ*mJY"*�E:GB�:Xk�������Y�l���2P1��B���1�u�),f�Va��VF��l��!����(�/�(�_Ԉ���������LPT�n�j�p7�������Q.#�|��!<�yUF�ߊ�W,J����, �
ipG��N�m���<���*ʎbl��g���فG��.�,(���8>X�$p��/"A�و�TFX_4^�Vp A���Iu��ױ����v\<�Ʊ�f��1�U'v�/dnQm�MDG6��� ?���&�s�G"�����s�R����笧�������i�ԓ��� ���,�S�Dh/c�V�rvm��1�Ƈ�(��/�oR�H����>UA���f^�)���i�if�j!���܁�~���� -ill:�W9O�1�f�F� ]ƺZ��O:�Az�O�>�^�\B"a>G�����O�!�_���o�j�!{m0���!Շ��ﻍ���V3�r���IYP	��B�ïlv�*� ��2\t�D��rT���o��?T��1��D�kc}�,˯�s�_�^��Γ����%�d2��Մ�>�
�=Y=�������[x+".<I[��dn���U�=ފ���X�Mi�ī���fӖ&�����˖Gxk3���s͇�I3��ѝ�R�l�܄r��=�&|udP�hr`,���z���%e���m�SG�]h��ҤZb5����rOG��N��T�s�H'VÍ�|'~&�0�tz�x�'\���~o�t�v�I�O�L(��f:��7eM�g:̈́8�;��ź�#��&��X�Qk����"~^�Æ������\����1�%���d��MkZJU�Nk5�?�Mrju�uc��G�n���~TMZX���{�=u��ǔ�bqg�qj�CL�kMҶ�^�j������W�m�*p�����\����-t���(�F��g�H)Ka*d�&*�E�`�;?uc���j`����tw���[=l�
�j_��������P�=�\�_��4��^
"@g��>�@_e1�2�}���!$m��~G��T%�v��9c���;ל�,D�?��W?����=������ę?���6=@���y ��bkUy�*���J-���!��/5�5�n�-:w�47{�V71��(5�#������G�(��ܡ&�}}�����i�{��5z��+' �z7nE
Q@��((\ ](W�4ퟐE{�� �ڔ���@�ڭm���#�Z(� ��E�����+,���4�@�v7��Q���mPs�V�$f���e��p��Ch@D�_ y��Ɨs��~�E'=I�%PX~��{��0v���+���*Yj�5� v�p����z�[w��5_j�S52�q��U������?��?b��i�|.�bj�k���.���7=V��%�T2�����s��(���T�-�-�-Dv�I�%�鮊S�':�3U�vV��2tmtl{ˡ64j��"=�[�����n` ����ֈ(�ߟ@{�:¥�l�*����5 `�%'p��S�C��<`��]Hm�a��еݬ��Җ�4���s��_\�B�P�!��YT'滧	t���Ohmכ��&x�G���kB��A�)�g�PP�!��<>���P*QZDc������S�'��U:�3��u-��ԝ%^X�#��-�VY6�J^�A{�'�!�z��������S�;+��(�'P����m3��if� r�|�m] �VT�,=��	�(k�������|z���ʁ䅰wؾs��3���v�R�%��U.g�Z�Pn!A=h��zt�t@dY��::�xڱG�%n�Ga-�t��^���(]��ˆ'���]��2�6��(�I'@�fӐ�i�k��X��PZ{jw*��Y+�}�nZ���#}RU�Ѵ�o]M�M�g�Y�*�nB '�ÿE�Qf�yu��W�B� �l�c��예�aЈ\���L0���a��m����~M F�[Cm=��wR�󰜅�,w9����|H�?6q����߿;6'�U�}6k��?��S�o�Vv�=��?�2!��f���
�kz܊��;���$y$ ��1	����%�ɜ��4��D��'"� ��(>Q1��`�������9�����P��m�o�fQC��Ύ�A�X\�w|�J���Dk�0�b��ג�݈���ל��uX��l]lQ�)�Ka��Z(0D�8������T(JA�~y}"T��rt5��	�]�¦��8�.�;@���Á d�A���(<�7�|�bI�yBS��荷ۑ�ѝH] ������m�	���p�$E�#��e���Z����<��ћ:S�p�R��ώw,$�����mj�?��wUP	�^ p2�c�H28[���� �#ޙ������8�XBH��+�O��W)�*϶'�a�]�����Yq�u��2ǲ&�Vqf� 
�K�갶u��O��e9��������n֑�Q���K���c+�}���'�"���Y��X����� �
����\r�����{���A���=QK��x;��E�+�&�b�C��m"(+ >\Z�q?��s��ҊE������tj`+8��/:�c
��,�''���V��,�Z �&_'-����Y[h�Pu��ZSH
9�W�b��� T�G�#����z��B��{{����^e�*tE�}�{F>w�k�_>�����K��G�+�r��R�`&�������4�fqǣ��!��7�s���R"4������F�����SJ(���X�H�G��"ho�.���B��r����.4��7k`����16�6O����\C��dWm_0@jlF^9�;r� p��
/� \)b#�
/]N�%��p�E(�������*@�5{�C��@�
f�ř�N$h���r������}׿;�X$�6�)-�Ǵ�k��|���z�:�-�݇�`t�H�E��@BY�����'�z^n�|V�������Ѣq��o���_����7�ww�m�ch��<W�8�r`?篁��A�\�v�O ��?�?�-q�%��i�nԗ�aّZ� ��ͯRs^�_�LD�$" m��N�HGFXH����Y��A�q�a��G�x(v���[���Y��"Db�&���0���D)��=VF�Ȗ�3:č����X���Yn����o�.�63ʏ�Ͼ8��Ѿ.̣��(�����PN���]y",=![ļ��g��~w�_������R2����7x ��4��D���3�B
�HGnHUz����_&|F.l�pzFvn�'}wm���S�ĩ����N$�c��M�B���W/+; �Z="���aС����b��-�����F����t�~d��g��.�LS�O�I�}@���{���O�ge0������@e ^�p��#�4U�0
n��o�%�Ŭ��y�t�zZvU=G_$��~����`�n��P:�L���Fr�De�Dj m� ��0�	 x��x�F(1N�I{��X"�Ѥ �:�Y����"�<I�I�
���q��i�z���h�m�{��pq�[����9S�x�z�SD� ��H�X�~J�BL�y�`[�N&����Ŗ"�7d���4�W0�Ή���6�i{����O��a��Z�����%l�d��r7��o>�!�!���B!�@A8�# �0xPW����b�2Β��lA\
*����)TD�B�Ó��J������@��6��pʟ��g��/O*;��C�^"{Y����$�*���G��.!&��?��ڳlrx����M~>��3�8
���CL �G�g=3���M�p��8�C����F�1{l2b3O���S5����`T���D?lw]�p��LӞ���l�Q<{����KZy�h+�O2����m��2�����d��߷�D�3(�����B��Fy�M���V�lIglC� .:@�nK���dKˋ5ا���``�h̅߶�� ��?��Rw_")ݪ���5�)e2�DG��!�V���6�2.�Һ�MJyy�ء[d&�e�e��b���{�0�r����9"3x�ڧhJ˗�e�~��R�w�onMCG�����2�΅v��A�(��)F�� ���`� �݇�ŷ����p���Ƈח��h(��³ʳ�{���ӵ&�Z3��޾�K�hv²�D�˷ln�:��N�D�<�*�������)&��1��flg��z��C�(2�w�Yx:q�t|���gA�HYV�)�Kۖ��==�̉zg=��s�����x��va{쭄m	��;L3Pe����řo��� �E�ٱfZ�����>�wV��5߷��G:��ʲ?t�z�ݷE��G(��3s��Z�,�[�oZq޶c��({��B��n����L9@�?d�9����ǑK��3 ���@��z��9u1����`�.�e�����C�+�
�# 3�#���x��yq��{�Sխ\����c�޷�=��� w�2�p��E��Dd�Y�b�9׭پ;�1�����e��Qfaq�M��o:8�=�F��	Q�u|�=k�������8����m�������`Zئ��q��vW�&ɻA��6�M/������AC�Z��D�������k���FӼtlx��N~�;<q���$3"}���V��.sY����y�j�*Σ(f1�2�P?B����� �nI�ȝk�M��>�`�)�c����f����iA��I`(	�
��� ��]���%��b�^�nI��x�׋ȍ^ ��:+�3S�ř��c���q��c����{#�eXY����:�B3Qs�7ZC^����B��9�BhA��ق�p���]��Y�L�jv]�(�F���l�Z�]�R�%~P�]Hs��m�n�����r��eI�ؽ���=�:g��U�R��_��7A[ ]��ʸw�f���ι�R�(�1H�2��n�*���V�N�-I��HZJ��P_\_�@�B��V�tАIdˆ9s�ʕ���j��c̃J�����@���H��G�e|v��������=Z�=һ�ir�-q��B>�ŗ�G��F�$�W1���/gX]|p�h{�?j��4DF,�0�H���q�'�=�m6s����K��b��#�w�2�O��;�	L�w��Lu�ˉ���̛�� �<Ry~!?(���0��$@