���6ѵr�l��~����I=���Ck��ؽ\�Y�N<$����9s��a��)�`C1]���of0uX����l��&i&�)�_jp4��tmk�K���`j��s�,V������o�x�&t�e�v���o�$jଖ�<��IK}}���h�8���n�[�d��J�?��`�.>&�r�KA!�WS�O6�-�1š_�٫y� CI9N�%�߳�]�6��y�~�����3�a�"b ��R�tL�׫�z2T�1;L���""�ј�2He������f�NK��&W�m}�}��R������E�������R������ӹY��o��O�7M�5�����r��ܱ f����=�Po�9�����g��w���Xn��G��c��3��^�q���U���)�}�TB���=���ܶ��F��}�:�����m��T���tڸ��ٮ^�v���9C���Me�|��.��W��w#���o�ym��<�$	b��Y�w��p�т��Ѹ�&�q]��7~�S�6�}yٖ��"�w���M`'Ğ���]+�P�'�\��t�D�A�� ����ӄC��|8q�p��5�lKOC|f�=�K}�q�E���m�D�>�p��aw�F<M0�{�&�����A���Kk̊�j��ֶ�`�q/L0�b�Ѽđ��-xPb�|iˎi�mq�� �253��V/����<��a��ȡu�>���l�=�w������X��^|��J� I��/�?�c|�����r����Сh�Gܪ0\􆛁`��tO��+\
���A����&�	�X�h}���/ӶV(K�^�Ѷ��8:n�J���U�
S�ڨ�[f���3c�j:�z��)KIv\z��z|���w��'K�_s��:B��{��[aA��Pb-�a�M#�VB�T�8 ��|o�<��P���c�V�����b�z�m��~A^#��p�'R�����8 �+�$Sșj��A��2��숰l����D%����]��ygf2�̧�ψ����BV��ɓ����8n�׬�l���l:�����V�)u[Bq|���qC�5!m���3c\֬�(�����ɮ���|#nCB���I����Ή������/d����盲Wh��Bgpm�0�]�[�;���Ǣ͢�\��m��Dϣ���}OT��*��̤x�TN]i%�2�k�V��V�ͼo�R�yC��^A_��)F�CUÖ�J�r�-��Ռ�iچY�z���M=�&���M�n3_��٪���)r�p�1����?/خ�����FBmȵ������w�o�o�_�ް��D7h�`y��{XA$WH��&����{�ѷ�yjo:���CcF�*]z:$��aE�$u�_��w����^JRI|��Gg���	Jǈo������g�ٽbfT��c�6
��d]R�y|��*�BՒ�����X�4<�a���3��Ӝ0�����Wu3�-��9����8�jM{�����@�t�)_�Gj����u�j��UZ>B��$�y�yI���Sv�MBw%�K�,M��BZ&/�p7���skR/_�5�F�t>E#��6���=�= ��>�9�2��-���/�ҮtY����:���Z3�ǻ�����|�q�k��ޔ$�����B��t۴�!�Z���`$]*<d��I(�4%RoRrs�������SOǆҾ��
�R*,��i�%Wo欼��ԑ����8�d�k��C�Q��.ݮq�խ:u̹l�V�Xc1rѾFݜC�����ԫ��<�x��/�-K����L˦u���(Im�ŵ��]�{'{�m>�a�Il��t`oޓ��yhqP~i���Q�5��%�It�f��$�J�J�K|-`�1!6��ȥ��6/XN�$�+�t�Ȫ��V����K%6�6�n�6n�l*�J�<S��}����YjT��4aF��G��fxO��164�Q��i�Py��-`:����ų(����$����;�󴆿�6�Z�vE���f�Y�9���Gȝ�=������ˡ��C?s�S �"�!b��>VTJ��d�%�����������
M�?'�Œ�E,`���w�z	rSG�ڝɻ"��6�]�>��Cɢ�7��'�'�DBZ���/l/j�|���a��5W+����;�S�����J3�M�<0պ1�2m����F����_��R����	5�AҦ���^�]I?�[s�#�!+]�j*�lz�{j[�l�H�@+G,�[���g#S�)�o$*�e���
�����	���0E�B�	��~�K)4%"�<��ʮ�~���y��I��������)
����9.N����e2m-+���)>~��-�T!�2�v���y�}a~w���!�����z�"�T��i�{ՉlQڢ��#1,�X.�(ըD�ڤ����	<���E;��>�=�bJ���1�Cr��e����lu��L+4L6�wga��X>i�������� ��c�S�Fp��d��wT�w��V�_`�.���H�A������ߐm��`���?a� T���@T=d�Q���5/��#�3�Ag�R���e�����]>9�)%��/��J�L�9��QY�hU�ݪx-�6�r�TĜ�4�S+NnE3ը�V�P�a�cH����Z]¦ߦ�N5���,�Q%��4��� ��uPJh\b��/ܰ�k莀���B�2��7�'�Yٳ�:Vk�W�'�������v�@�>���hp��,������d�"$L����C{�_�%�����%��KmLmX4$�M����C���$�M�s�%�������x�����SV<�N!z�¸�a��Ϫ�+�[�x�c]��&��0��&�"~���Հ�1��0E���������9�;��ن�&���?��G�&Y�������;�?�;��_x�X�&�g e3���m�>`$hUx����Z)1lL��%ڥ����ʦ
���H�5�X�LIc�\�	W������l˙8[
�C�ƒ���u��	���w��ÝS8��[R/��X�(6.d�t��[�Lᕬ��<���h+�Vn�,s�c�@s�|���[D�g�Й����T�HT��O$UV�Y5�j����O�������9����]��ڂ��b�
����������	��}��}RwX��F��?�4�qwo��a�����G�G��>�s�>`���=���cZm_�@8�v*Ԋ)D�}!5�%w�`_��㧺M�:X%�Bd \Y�'A��������ʏ|A�2��F�NMO�~�v�u`g�oQ���G�kAƧ�W�~Y��׺}ںi{ۤW��L#��i�s��ƨ��w�b�=qk|�ωUkvw���o O_�P/h-{�w�.:ĥ��3+��1�>���GF�?�+���h�L4mxȨX�M*fQ�B��<65�ꃰ�uU�|1�?�k�t~1좨��n^����e@LgZie�ŕuh��A�'��ԱB��F�I���E�W~U�Y�}�~�w�~�w6x����.mL�1���6�j�5Ѐ��[Ֆlvi��>g��ik��;k�^ng��af>�7q[�`�,N+"*���p4�z�Ah�NG��>y���5�f?ҝ���uq����*X�~��wͶB��z@�j�'kش���5�lc�:P���RW2>���B�2ٲX�B�2�U��L��}��E�o�#t*��@���SV6%ʘ~��̽˲C�6�m�Ʊ�[����$l	��I�
�J>�l��l���J�_��I�t��M�O��d8Re0eB$����Ȥ�cZT2S�f��h�?���f��I�bY��
�:��`���2	C��K�f��p��X�̍r^���`�}�y��N�Jb[����ܹ�X9"6�	F�X�A|5p�9K���V���(]��.�:�Ќc����*yF�=�n�tπ5K֌jӌ5{\���(԰v���*M��rd�a��nU��1�*L���U�CC�lQ� �d�D�D�D	8uI�
b���$�sE���xXày�H�u6@:���p?㬍�p��~�mmr��	+���U�:mX5�n6.u`Yn��8'^K�30q���w	�����o��i�G�K��v�^�Qb�`�H
*�x(��@H���K�A&G�tŚy�J�s��;4��|et���&�wk 6�a:}&��\��N`i2�EL��T̀Q�
.(�Mug���t3"�r 4�cS�`6�W�l�sLF	
P0#�o�y5��̀nfeH�B�v��j��be@������M��M���&V$)�'ezՊUN+U-�d� �{1h�U{4�҄2+͠�H�:���Xs^M�k�v������v�Uϖ=bu�e�oW9�
=��|�d����d��4@RUl��o��1p�7E��=���
p\6�h&��������`c3x�Kb&ɨv��pXoZ������g��C����	@�h��Ż�gXL�-@���n�!�G�F��&�֫�Z˭M��m[��a���'qj!Z��hɭ͠i��g���נ�,�8 xº5��h��ot�˵��7tP1D�' ��1��(��L#=�Q֨Z��:�a ӥ�� �W�?���סw��9�Pa���W�V[�x�U)`�B�T����h�[��}/�
��9׫@_��pBM���T\Ҥ�+��`��dX"V��2�wZO^ߟ�K��%�9����ATÕ�	��o��;������o�o��A7��Y�
���[����k�c��<O�}�7����A�,��/т	�	"��Z����1n�N]`��2Ǥ-2�?�o]��^޴��٭��]��l��]���SR��Cݴ��H񂯐U��G���S�"���Ԡ��Q�����\&������~_A��u���LD�����[�:�X�\����׫��_CS�}n�����W�v4NW��W�=��p�(�ݰ�_���Ț{�K����#uv�+�x�n�������z@7N���_����o�(<��lG��,�R�����U�+p���8��@��_(�9|��Y�z��K��[���9~�ꛇ���s�ϱi��>��z旁���A'�B��4n�_`/��H������?�֜�i���@�-�W@ɲ/�~��;З���?�zצNK�����뭴�ꮛ��(Z�B��O��9S(	�$=1��P+;n�0�dq����b����z���U�v�BJ�dA��<}�&��4`�{��g�����f��+�,���c��D�!�,N����}6S<f�s��{�k�����R3+�ƟE��^�]��' nC����4yƴ�k}��$���ò��� �J�om�׃3�G�����2���r�s��=N�~-�n�1� �VK)t>;`',��^A�תH��,���m�t�\*�sxs���H�X�����b��Y��9A�͝'v��(;C���<U�Q.<2�^n��a�-�&�^i����=���%��tD��z�tg=�P�g�C�V�5WJ6�C���;�N�g�5+M��^�ԷK����)�c*�)$¿|�]�1`z��b��W�J��S��B&q/����b '[\��P2�j&<�!���u��@�l���
��
=:ts��V���+������
t�đX�!!)C,�F_�X���<��N�.�;��9�f��kY�"�&�5�M@�S��|���m���;��[���7`�p��N�����B����ypPq�PZ����K��B� �QgЁGy�,�w��{n��e9�s�e�˱yՁ�G糧��	�#[l��e,w @2�Z�>CJɼ�d�H���t�L^���M���
.�ԅ�('b��;s�,��lZ7�;_u7��5���N;Z>C�jUl�z�W�	��#�o�Q}4�B��c��cC'�y�t6t�cA���o�a�f�]���$hc���%.Ug�W��P��v�yhQ?�2�˞J�6��=����E:�/E�]�vĮ;��F/���й�v^n�0@��Od���CI�R+���x����9�B2������v����m�9��F�[G�4�x���S��뭄�c���b
�9�{TL���t۠��7>P5D��=i
p�t9&�����Ȉn��Ԝ��$���{| ^�.�W�'�k��E���<��ۀ���i)�:
�{_�;ص�A��my<��k�K�� a����N��P T�F ������2I>� ��SL8��D��Vi�!�z��@�3A���!�V�p��z�i?��	���]H����&�v|���!��tä�<迎
լ��������3"g�ktytT�M�r@�mİ�ha/.����BV�g�5R��rqBr��*Zn:B�64�?�bs����e��<ɥE�d}l�$��_:�0�"z#��y����k�uh ��T���7L&�lj+b3h6�46�9E�ᗳ��6+��.�EbΞkm@EXh:j��1G'P��_UX����}�M��IY.{�����ߙ��#�Ű���0�B�����8����|Y�|�i�UR�� �<E���(+�k�P��ؐ�}k�����4���ޡϪp
����p���C�G\P��G�nno/��[!~�0��W��v}���)XG���vQ�>L�p�. ^wHBF��n��ܢ6�jv���JB�oN�8#�j����*�-�V���r��4�f�_�X<��"?.����p+��̟��㾋��8�^`�-9u�,��O�$��6�;��Ě�y��3���8����M�?�y�_���B20��(��Bu��w�Xy	3ޣ(��)i儺��R)h�H;DƓ2�5��$�$E ��&��@y��|���#������J���Cpޯ��x�%M�	���/43��ǰ��[��h�g��,�EF:�5ݰw��ۋ�:��]�l)��)�OMJ���9�/غ�A�m9"X3r)p`+�k���������o�eT?�) ꛓ "���aea���6^�O���x�i��z�_�ՐP� �^T<��0��y�8���$�ٰ���i:�;g��]CE����WY�x	j�>�TJ��g�jC���/��º�#5b�t�|���]m�y	d��#r���W��aܟ��U�HjB�����Iۑ.<	���W�Z���"|8�n�%�$G��W�
�g�a�N"WHX<�r�UK	^R!�����v%Ե��&�B����MT����;�F�Z��!���ޓA_�l$�hH׆ޕ��e|��	J�褙��jzk�;�oo���T^$1�"@f�L���� �cc�3Q�t^�exNg9�^ۧfFgO�Kl4^K&qjD)D��ROl�¹�x[��k��<>Q����D}9�(LހLkWS9�U>�5���&�2����Z�bL<x.���$æ� ����/g�&`�&��iŦ��(]�g��Ϭc%�!�I�����
%t8��!M�j�EZd&S2�c2,��3yhbe�ub�at�'i�k��슾\�� �<D=�kUD;�i>o�E���^F�L��ai!���#	��}�^����܆u����)��8�:00lۆ������3��A***���v���㧘�ag���c�>�P0ϙ|�YXDޭ�� ő��r�f���e{)��4����9�w���9��Y��ٮ]Ԙt�k\����P��L����8��~�7�`�!�կ�(˞����V-����%�S�������S�I"3�N{ ˩���Kz��G��4T��� K��H�����O�d�-�>w�T����k�ʩY�ƌܐ	��1�U$хI�.uHi�����[� q�A��]&yG�N�ۆ�0b��̒޳�w���ݛ��Gi �/Y<� ���.�����"�����=�㮑h�&�hl�Q�R�
-�,$�3hl�P�>�V���Ѧ��2(�����q�j��)���!K�0�u�!������8]Qo|R�`^��XQ��)�t���Y��#ƛy)���~��y�ZOw�|��F�y&q�kP�[�]+n{3%�	�l��x����T�LJ��!{���-*(�ˑ���j�O��;�z������]��#���.so�=��x�C"n~P�8�t�������!��a��&�j4�Q�@��#1sJa��Hl�;��7V͕�����;��k�W�RW����w�ws���fk��oOZ�K�Ŕ����(��q�%	�$�f؟W򣓼ߕ����C�9�
V�\I�]�Q̿$�Ӆ�R�d ���5��o�ya��eC������)M}����
�LDm`A=¼�}m�Dk�v�$���gM���q�򞺩<��P�8�̆�$֧����ȕHʝ��n��< ���`�ޯ�+My�0Ӟ�_*\�I�n(-�t8~Y��-|��	�)|�6�9T3�J-�Jʧ,?~\ⓝO��2�[=�L p�3���
���A���3���!����צ��l���&�kY�-(�̊��T̴���O��[k�[M�_ ��C�F'�^SU�X 
�,w�e�Û�Gw��܂�c,���}n6D}��.�gbp��몃��l��@��&}ͧ|���!�����Ca]�^k��<Ź ��<@�<�Pd���M�4�=F2�Y+��ǵE�(�k�%ml%[{PRFir�-�������tir�U�$���V�����ҝ��qoO�Ÿq���uk�����UO��L��������,x�{����[p7�X'���S�X�(�����kaO��ʉ����C�b����k̡Q���V�B�ŻqU���^�gK��`�ʕ	�rHq���AGOh����D�yhۻ���|4��:��vנ���t����+�xuT?�<[UTZ��ix*�QG��P���3�㗸{����AA�i����$�Je:�����}��"M���`�Q�c�eRt{�����W��%v�]�U\�5-mӐ��$��'��:b�iϪ�ud�:���,(o�r_�c�oUu(�$�cC�B��*bM��},V�dN��QO&�;}Y�6w�.�
Y���� �W&e�@;���r��B����6���/Iz0�i4x�1�u@�m3�������6|x���Y�mP���?�p�N�=��~�����2�z8T�@W۳J2��q���>�X�l.Y�����:Ɠ�����ʏW���[>EU�]5���oH7H4���>�r�m=^�\�dLַ�F���f��o۰��h���m{(&��>Kġآtm�F����58��p\�g�c����Y��;���{P\��lǾ��W�x���]����!����;#!�U\ןѳ��L�o@%��ӿ�՚���U(ZvT��w9�s�Ѻ*N������Akm���|M�b����ct���
ou�)�$��'��<r���Ux�x����8�σ�Ig��}�����4�9 R���Tԕ���&7����Hv����T�b�H��`3@ea-�q��_L`wc�A���-m�9�tc�ƿ�����Ϧ�����en(�ѿ5O��u,m�Y�QbWՎTQp����IğQ�ˌ�J����:��Ga^,waqԓ��e�Ȟ ��v�Vv	Ε�����4�J����G�t���`�G9��*���|i��2GA��I�` !���S��5�8��� 6	z����bChд\�4X�~*�\��X�ς�%�R�Ԧ�a]IM���j�,ݠ��,�į�]����j�k��="h�j��ڰ	�`ġR/��i��Ĥ��%������ח�\m�z�В�Ɣ�S��c``	�a�qD�[���;0�C~�_?��vp�h�Q�S^���):���nC�tz����ѯ9���MFylz����@k�Q+�N�r������8�u�3��T�q��'��[�a�\�P�yR�>��]�Q��&j��}U��g_Se��H�h  ��0�}�ʓv�]���O�����=�7�t����I��>�O��Q���+MGc�)�4瞿���XԶ�&�|���<AvI���������9~*��8<Nr�|
j9~]H�꣢�P�Md�IBk�At����WO�^Qm�w��K+�7��,6`o�����E��*`o_���Ï����=�̩�R��s�T�uHD�%d��^5��΅���n�V-��j�Rk��|�nw%k��1��LK;�S:�/urt�P���t���B����x?�`����� Fe����P��;J�f��"�Q<�m
^���ϠrM	Ed�`(�q�����(���W�t�u��������I�����ԳG5��5%�5N|:VoT�Ճ�t2/�iW�J�"��w�YZ�G�!7X�S^U^��7��~��f���"X>�^aP���X�H?v3��J�f~	��e��lO Չ@Dm�R1�]t֔`~7J%D�mn�"<;�6, �	�`�Fݢ�ݹR��B2����n�x,F��{x_��?��/A�</���lk.~~QT%�Iܼ��$^�l#����z�������&DxW�i
�n���׮ j����� ��K�Â�d����F� j殭&-e��(�4�PQ����g��N���P�p���P���"S7��Qq�=zE ��u>v$�����9h��hzec�t
�yY����m^Z|��K�}l�xd��U<��&U�����N�:�/TDu���.���t]��t]�S/"K �q��K�
%������[ݥ�}P|���ςi<*�6�U|+��)���U|�w�ag�d�QL*>xl��t!��I*>,).��J�����]��+�������F�v�C�+���S��&#7���*؎��'�طZ'��:>��㛉:9�Q'��3�kh�M�}�I�*�.M�6,A�yai	���)��>�#�a8crj���������f/�J��a%�؎_��O�4/�J��i���7k�pyM�kx��:��nK�5%���έ���}���P���ŀ����VR�HS��4�R���Rۋ��%���^�q��[��R��g���}5��JpU�4��B�
��!���@�Wj��x����H]�ȸ�v��m	T$�xYӾY��}CM[o0��48�b�L֝9�,����Z�S�k�&�s���'��nU�T��I(Mb{*d�+wU+�"�wWW��77�I$�Z�wwq%�ηT�� ��Q��Qm�q���C�HVD8kaw1l1��[��ay?���(�.��1�	��z\'6EP�r���[�;.1�������R�cF�W�<�֓b�`��F[�A��Ģ .�b�j�w��,��`�[=g�V�#vx��
c�TS�gP +�s{��rBɨ넗��3Q4������~o5wd#�IYv	�6�XN���E~�l��{��Y��a�b�h�}��Բ�+l�|�C�ꢔ�JܒնL�N��K1D����/��Q��6X#�y^���!(D])��x-��r�T��J�}������k�����Ϧ:9�&1�j�����߂�S�3� �Q�ϖ>B�$C��6�`��.�t^�z�5h^Q���mt��톀�2
�G�_\e}�������W��i�$i�o`�Hy��]K��
�g�m���$��S���
Oነ	��G+�����T!���-X��,R�tϥ���Wp�����>Vx7v�̷Ƈ��1��$��IhA>��/��P����˿�q}�����;��N�z_�7?�#��l�yy��,�D�K�S;>�?�V����~�����[�b���kU|�"�U�.	���T'�tW�]c�.�{�Q�6�F:������U�f�! P���F�s�^�@���u]/��#/�Q��
v�"bTxbpe���S�W�����z�`�E2/ceCmx^���_������7@h�)�V�y�k�=��eDy@6�k�%�C�E���/aN������r ��f��~@#�9b�U
a�[�5^U�S��r���ɩYM	4TC�ѶŤKţ+"G�\�vrO�|L�u��Yu�h[~z�A�RA�/��D~7(���+�Ž���Ά�*֔��Y��d��V��ʊ�X��e��	R�l�rY��,ևGE�g�����I2R���b�h=V5�#MV��%�P�ҁ(�4�Qj�+��E�8L7(5�@mUzzX~��Z;\�����Fq��r4��1R�m�vf^�z�)��=�dÀ��Ӎlb�JU�/A3�%���� �z+��|����ԦяA���8�qn��O(C���s��"S���+�X>�f. U�_��$�y��u�><��Jq�I�mG�UI���X��ʰ��	������!4SY�U�EreRY��q T��J��]Y�eo�{1>M�X�x-4	jL��o+iS��\�����%�t�^G�6��񊚍���*@�~w>��eE�C��$���V���!<��t� ��f��[��3�<Ԗ_9�5OEU��{�0h�9�qn|"��yn|�F��0�L ,���j�\��̱��A�P��oԩmx�Cw��Xa��N(�3+�ũ&U쀋/a: �K��\�����k��I;�
BX�UB�x�WVP鉬)��->=��^��Yp�֓�|��/��єc;L��� 4
ȗ���טC �����Cj+p�gV��R3�c��5Չ��Y`^�8zk�RO6D��)��9fZ�:W����,n=CJ�y�$D���p���MF�5��v��瑋��V&m)�2'^9'�5���Q������#J���q�W��9i!��'�Q�� N��G�s�TyJ���7�`��8��${k�s�:Z}!T�⿚��'p�5�M��L/�? �4��p� :��eˡ��5~փ.�f:'4V�Y��c*�\��U9���(�*B����X�GWw� {@e�t�ˊ���*А�%���C������l��Y	�a��r�b\K�+(q%�<��*E��|x�fÿ^90��]�~�N9"y� �J�R*��oo��O������h�=�T,w�8�U��|�H��7�[��}v1:�Z�QD	(}�	�_�0������l9@:��켃�u�e�x����i,B�K̡�����g�������#/�͉^,F�J�,��;�Ɖ��"6 �Z�8���vd��[ot"�Z:q=,s�~�L�U��V�gX�
���S���:�6O,<|J�zV��/�b=b�ҥ0��}qh��s�\Q��
a���&�Ԑ��%�*1��#}�/v2��.:Oxq����[U�{Z��w*�y�$>�ZS6�LCXaEu�<].���KL�N�=���+ʕ���݀�����G���	B�y����`�/����U7��v�G*�Bh�чỶ�e��ڏ�צ"���h'��W�<��V����������^�
���co��'�djp\�@eo,g��Uz�WH(`�������D��x��Pk�8I\z�F5��x��5�}��C�S��p����ҿT��`��Q�0���맄�i�ӢF�<%��4���}�.o
D��OY����p"�1?]�i�\VG�zȚ]x�7[��Z+�w`]��dh>�����y�$���2�,�r���C�o�5n4�kg�FQLQMZ��<�\n�r�jFw��-��1��"tqEhjEEh����%�݅]o���]�ON�k�'��u����Î����Ja���/�M���l�G=&/��'a�hV�uÞ;��6�����m��ȭ4()��2��_�7���(Y��Ü&À��A3[pW�mU ��KP>P=w�>A!�����~�ĸ;j�N�:�u�v�`�i}h������V<��젱�߈?E������Q����3��l��g;�au��A��/+������3C��N�b��P3�1Z)V�:Q���Vh ��@�����E���jе���D��V�`�WzN��YRZ��̼q�H��1�DG�%JK��Ē\/+,E�&��P4�QZ��_������M5��N�A��RώT���؎a\�����]�3H��.V�b�郀���*i|���x)�V��d��}`i�2i�Sv������i�tV=��s�g�E�|%� q'ƛ9�×8m����ٽO�P�� E��� ���b�@�MoK�!��ai;� �e
z<���6����Kx��a���#�6ʙ���� ��|�d��){d	@�%�jI]ʅzj�~��~n(G3	�p�R��IS���Uor�2!�3d����H"ei{'��2�9��]��D}��J4�T2�U�>A#$:zx�����%P�xo�|��"<���ڲ�Ӗ��-nĴ� �? d�À5���=�}�0�+H�L� �i~7�s�IMWV��3R��@��
��υ����E�Y�0E+�Uؑ�m.�< r�ʋ�rl@��5@6,�mX�혥�h����'���΅�u���R��4�e!��n�h�<��3=ќI������r�U&�<��0~�\�+������-j�:��a;fzFE%i}{���th�i4B��bnʛ�C��O�8��<x]��w���-K-���1c� -\x�%8�A\e�Mْ�`q�[�1[�㜼�D��+�4NG��/� �m�,=p��^�� ��*��-Q-B>G �����)��+O���!�f����g����G͒�?��QC��Wr�X8��oE�ev�ߠ����,�c`�[�L������Dn�_��E��d��ZD��zA+�V��B�a��
���؎t:���a�deBn^/w�4�ݞ���8�ѵ����"�鱭~��Q����*��7� Ix�q1��������<�{����-=t�a(�ݡe۱V��n��{v��t=���s���P���#�B�gi���.�Yqe��Ȟ ν�������6��r,]��d);u9G�7�9x	T�;L�eco�G��W�O6��c���/T*OX:sDǡP�����o�ǲ������ݏ-�p�2�҈�:��p�fCS�%+�C�	�R���5��0+Z��r2qV����J85C͹JLf����2G%L��h:��?�n����V�%b�u���6�ƅƏ+m��M3y���~�X�`D7�5{S T~�:;ov������_C����`���:��N����p�	��dh��E����b�×���O9�
jk��x┳��'K��b���)��Y�S r�il�܊��2V陃�+H*
�9�4��Ԅ�c�K�3����MR� �~��C�x���-���N9�z�P��4�������)a�V�mO׀��"�c���������̞���ܑ�=SnJz:��h�'�f8��	�R���5Ҽ.o��aM�nm(�$
��h�%���[�\�/'l��t7k����P�4�i��8MM��� "��!��B!q�
3���:��v�I�\�#m8�l�;�d�������5�Ӟ
gK� ���=v��2�g2rM�R�k"�;�5�SA/������D?{���\����#����>�Xۑt������Ο�t����X��l�+��%� �i������E�k��ז�m���(�Ue9��D��	�'���u�uG�w��r���,m�zk�o?�*�)�ܢ,+P�k�;\��P���w�d��}����g��T��� y25�^���NDƫ��4Ր�,�~XY�'�ށ���l0���Cs���I,��-m��
`��uv{*4��3�ԍ�c�(W��zwĤ��>�����t�*����h��v���}ڟ���2� 2��6�3�o!��n`Q *{��|CȦ��!|1pi�X����g��cdkRO~Ȍ�|�=�_�� �^F�$�%m�������� �< ���c1�Pi���f�x��%�Dٺ�q.4� bگA�\�8,��@G�L.�<��E([z�c�ȅ��s�����>Fo�QABnb��eI��T���O��؋E��Ф ����3ۢ!4�Y����xo������TPK��(��5�k��Q�Q��l�f\
�K1w@ms��g}�h�´���<��a��� ,/OzO����31f���b��|��O��+X�+���c6Z�Y�&ۓ���5�
=k@��<��Ҽ��ȋ-[:����K��c��hJJD�͵x�AR�#���J$ũ~����_���B�`}�g�`�#��Y�����;���No|y�~K�>d_~L�͏���'��mK��o;�ŷ�-mw�۶��l�w�x��W�#W�]`D�E<r������!g�@�tg=�8˴�}�&�<�P�1<��n(4
��h�Q�g�cY��[��ҕ��Vsx�ig.'|Q��&���%���@1��!���^6�Rt[͌�0غ�FY.��O��.Qc(
��Ygiܳ�C�&~�9a,�h�u�����1�e�aC�I�cp��v�/;�<�	J���0�HF��?��<x�B�����iK�C�H�L��-O�r��nwP�}Y&O_�nM�'�������ٕ8-��x�j:w�5D;zˈ��ⵓ5��(EǬ�2��uB�7�,����қ�k#��)�|����,�܇lȋ�wX�k�t��VO��f�~@�h)
 ���OIb2�)�٠�eu���!#��6,µ�J�L�e7�x���U����w��J�loZ٬B���$�^d-�$���m�~�ӫ%����!����Z�׷k �!��1���v��7��=Sh�B�?ӱ��39�xE ��z��z#Z.QR�S�3�8u���
c�Y1�c�+��V��41�fz��7�7��Ab��9�4� ��6�_ �����@���_��A8/�m�~�O��M=Ե� ������:@���@_���)E�@Y�|2��;|�>lf�)�z�� |�$�'��Q�"�83���t��*��1L=��!�W��RH�����:;����g)�E���
� gv�lǐ&��S�|�EJ;0q����?����)�����t�6�(3@(��KG���@����|�Nygl���d�/A�~����~R_@}r���u�	H��f��`2"<�X�_�>�ݺ$ދo>1�3�eo_�/Ý�p�^3�.F6�L�~^GC�^�q�;�`��5j�9R]�)��E�����Q�{&���H�F�����xR��A�}�Xc��?��h��1kUT����2��4 )ra�)�8'\�ӉZ�����ʓH�)NK���B�a��猵CT^�1"�*�dEz�r}9�0W%�Kq���ϱ㉋t��2i"|��i��]��������w9�+���g������ց�F��W�b Z�A���!h���n��	��`��. ho� nd�oE��o@�r}Ω^`�ѵ߾�de'���@��R��;�]x"�b���4(j��9�r��]/+v�UĞii�	��<,C#��2��W�����Ph��jȾ����ER��_�;y���>�?��]���IE�&�ڃ�J/e���?GE�+R�z֪��I��w��+�P���-��W��Ŭ�@ށ��E:J��a�����zfk�
.ͤA���lm�ȫg ��SU9Zk�y�r�_>��ger�d��N�I���өޱ��BM1ވ������GPjJ������0���>l�i��HS��Y�/�JhF�]�� �*�|)��_&"�4����s����'e��ja�^LBn��s����c[/�,�t�E۶���e��ɏ��*�Գ8�{v�i"��bg<q�[T�kQ!��)�;N,d�f��2��섥͎) \C��l�$S����3}Fe����kBc� M��1/>
yC0�3�r�$�5�)����6�(�!6�~�aA�Ӫ��٪�2 ˒,٨����vl3������o�Z@ce�g��r��Z�]*<�
�V���٪.x�+�+�f��D�8��� v`�V�Bh0j�[��+�!�t"��V��$g���S"��� ��s���
}�a�V��YFU����ay�m���#�0;�p�~`�IZ���G�m͒nE8�g��� ր]:����g�_��i�8CB�f��*[߄-��f���a��F�f�>Uk��P�j?ni�I����$�wq�{p�5�h��J̥p6Kڡ���4*��N�>A�9��7�J?Ы��;�2�. =��_P���F� �Ⱦ�NW+�z�mSP�,/s@1E�D��:k����)�(�Z�Pu�&S�8�)W�u�0?wZR�������������
X�df�x��ɰ�'}ڸ0%���J/p��ǥ��F��ÿo�O��_v���+���;ĎA�N�&5^>׹�x:qR"�h��AJnݭ�g�]�9��g�e�ܡ+nWb'чI�lR�����G:(����&h=��/K�3b�/���(��r�xӑ����2��4�B{�e��I$�`i�=3kJ�x���FD�G�q4���4BU�G6��3�K| vb5����E1�����"�UF�*dl�'��*}�o$�2��H���lr��z��ͩ�R\�)�pBO��2�q�4�K'Z���Ӏ7���d/���.<p<\|�1i�hZV{��� �Φ��L�ǝ�PIW�Z�;�pM�ӊ������h�\{���?��C9j����V�OC�`MӼUU�z�T#��M4t�45p*��O5�ï�3�E]�71�=�����i:i#M�ᵩ�;Q�Q@OZ�i*m"v�h@�ziE+��F�	�F�_*�
 `��i���r4Y�)�+�iҜ��.�0�8VL�����)x��JJ~��/v�K.���0�D�sJ@��`}~�1�4ĖN� �0XE�LI?C����K�b�-m?2k�P���=�Z���^�H�S����x�-5k"]�`	9m��te�F��z�����R�>Q���|Xi�dN>1"@$�5ϑd��Ҫ/�Ճٱ'P��k��������Pk.����}P�\��zm?�?��;��{���b��t.�}cJ�E��r�H��.�F��y�=̔�=� V'�x!��76Dε��'�'�^��F�HF�L^��ǋ�I/�6`��C��K#���N��s���=���K�:���<����T=�p��&S2`ˮ*(�c8Z<؎�W�������Fˎ�f �"V��6"���B���d���������/м���� �^��^z	��w>/k�@c�va����A��ɻc�#͍�V���+�ș��r��Pq���@%#ja�����My�YJo�)��YگV���Ѿ|/��D΄���a^kFW�6�هj��.��x��xCs���!6������o��/��K����Lb�����gC3��9_è��9F�0���yQ�p�<�)�]�@�Ԅ��g��	��^i�ޞ3��!V@�-C���A猺�#��DuN����O<�uN�4Gu] ��z/���X��m�['�i.j�[qF�݂Ԁ�}/��*��H>қj"�%���D$�����?�6?R9����Iw���h��;5y�h[�I5e!�
D�XÍ�N�����^�CI�]�����W��D������m��/��������YoKku��*;~@��JO�Kyfth�6�%��C쀠yM�OěNnJ�k���P�u?�w�ݨJ������Fbk#ݦ�&��T��{�a�"�ɵlۏ�uy��2��vM�5Z��M����vhF�M��nMx=�I���.��``��3��w�`x�����I�R9`:d�õ$�?<AM_T�T2�S9^���Ҕ�a�N�!}��$D`�R��2�	2虋�~������0���Y��>f���DIj0�2��gߺ�[ǫ��c����nm�*�I�?���`���ֽ���OC�PްR�;yΊ'ȵ#=��{�����v��4N,-R?-;��n�L����?t?�=�Ζ��ˣ�Ҵ&��J
��(b���̥}��R%�a��+�)OT���moӶ�إ�T���~?���@y��fkA8�TY�54]=f��=�AV6^��� F�{0����\a3(C*����^5k�T�|�A�{]���D|j�X�	�PjHq�P3%��E'�E�4��qzV��Ї��i�g}�$Hpϡ��ż>��e�ub�8B�� :� x�W�)g����5��l� ���^A��@b�Mb��)����5Ne<-m�(Ӈ*����h��/&�K�m�Ȳ�+�̣����h�TE�X�*Z���*���+rm�Z��|'?��;I��=h���-���'u�(���M�Ҡ5z�<{��P�������� HIt}�_���*��HҞD~��r�������w�~�@��Iia��W��3�:�ڂ*�Sh�;t�=��p��'�M ����oc�S̞ɕ�b����_�T��Zy��eG�P,�W�`ه;�u�a�7mw�S8��(��1m?0<�̑�d�D����0��;�@(���3L��̈�\bU8EPR�g��3I67F���S}3[��窬%]1�)�L�� �R�Z�n�p4Ϫ���$�H��&*;�b����f�_Q���^[z���;�R��q�Ϋ�Q��^*�:�ئT�b�:�oImBj�x�0a&W�߹u�Jp��&`Kٻ���,,�E;�&��q�����	�%#
OK�\Lkn���s�1`�G��ʾ����1� ��*�06!�nP�����9=z��q`��ҹ�!D�_ /���WZ;�4V�1�@<]���T'��h��p+>AM���0^b����w��c0��lMItik˳a\�g��?/F�p6����l_�ҳa<҈�q�/�\D�i�ÒZ8����{cЎmE䈩m;0k�b��.�YR�ދ݈��ˮl��Rd�,��	�7s�2�O>���m:z�V�x���e���I6��#"0"�l�=���L������i��.Eyˎ�LL���וNǒ���c,�n�ě���g�8�i(0$h�]j��Nk�ch���M���;qz��f��(��g��ѷ;�jHy�Y��9v�E<���o�6���,�p��Eϔuv*N�j���v���+�1[�E��}�4de
����k,)�Fe�p���_��W\�g��>�����&� ǘ��aw_&��%��19�&�����!����S�9�֑��m|?���%�� TƑUǴe9=�	�ޗ�l�L��O����X���Q�	J���>ճ3�G�97���+T��d�b�M)�U�EYV���{N�N�7�`�G���J����*�g����j3�	��p����k�Db�	6;K�K�K� ��7#�2�{��9y�U���"�&i�W��*�T�9\3��We=�ߌ��ВS�¥���6��[v��tl�G���&� �`ã���|"{w��X�#]��*�"�~N���h{}!wRف7�Q�5L)�"��z��.�O�赑��4�X�j�d/c��A"
���((�)��Jw����h^m��>B������y�"kZ�r��;��iT�^!j�Sol:��_��^m�����C�@-ܖ��)P7��v�I]}#�!&鋈��Q�U��[&�������EkU�V�I���ނQ�G��q��|o-�=۬$�.��OaLD������S�hi�,U��^��QcDwtb�K���#��<;��*���7�N��������0�Jit�^��aڂe�o�)+�qz�!u�H�825��5�aAj��*�J�lj�A�.Yv��>}��*��W�ͱw��&����o��8y>ǳy�K^Q;��82< g �HF�)ἥ�4���V͹ QM���������J�m8�C�TS���+�7C=�(�	ၼ֖E���Xv"�*��csAi.���3^��y�k)x�\���P�����l�$���.���xw���h}��(����+�*�����%�,?�Hi2CSTX�	����Klp&^kU�r3I15@#� SI�(�x�ׂZ<J:~��Z�$̖4s9k�D�1'rت�̀\��v�Iɱ�X�g�N�Q�n���x��]��^���ҫ�ª�����2{]"\n� t����]��M�V�(�6ith��4���H��)�-�U�[�q]�|�����k6B����G��F�u�`^����s��7��*P�-���`�6H��dKyb3h%�.:6��U�P�༉w�4t���,�R��#b�b�f#���
Ò��;/�tΌj^��^)cؽP+8�;�m��wA宽��Y񤞂]ح�ZP ��z���dEt�O��b�ޅ�����B�Y��	Z�E���?�C�0�g���X�c/=�[;�M�Q8�4�}9E]�t"���� z_I4gK�b�����1���b�Ӏ�o~�`Nx?��V�F�I�E#�KO��)6a8=�pMtK�1<%=�=�A5�A2nF//�"�D�W�0=<���7-2��+���nI��-�������xL������3`ؘ�i���T� K���vAw��\9PX��3	�[=��v���� �^5�!7W�����t�eM�;P%� ��L�\��F;������7�`z��&זbH)�!?�7bk��uهj_S�Tq߀���ꁷ��1�Z[O�+�M?H6|X�o\�8�L��ʒ�_���^W1�_g�r�'%bH�qK�K�q�W�����`���wU��u�i���y`i$U`��6Z>�C�4�p�P@�K|c(]���M�t!���Ǡ{�[4�Jy+F�u��y'8\� b.*B����O���$�
)<�*��V�^�e�z�q:��^O����� J�Sx�b���a1���|��44F���9jR��F=䯱\�H��L��|X�IL�����;΅'KϞ?f��Q��g����C�3?��m�,u��>��_J�'bLmʻ�?{�'`�ҭ_	�3jʒ�I��O������Q�2Q���Flh*,qx��d�/��'���/�U�����`�����z�v����p��v;(��:s�X�c��y���WYv�@�?T|R��&~\����\�Kz���p��7
��
PNF��A��O�[�*e�߄�F��xq>���:]�2I��t열1�*����K�K��z�8��������_+�u>@Ph�ỴN���i�<����)(c1�� 2�G�"W���W��Xh�H��!�D�X���2$nE�d�Jrӽf�:i�c����N�RD9��[��<=O-��FEc-m+ɶ��Hv�T��=�1�9��f'�
V�H
����2i7_���q@����*�3LD+L�~j�+Or��M���M�dSr���J�~��ݔ��dSK�_��a��g"cd?�Y��'�j�(	����1Z:�[:��><�a�����4�ʓ�w�|ܺ$7���sj�GL���:1���sjN�k�ʓx_*M��rp�C�c1�j`Z���L�|~���4��)cUl��M���}� ;�6�O��B�.�x>�|^�x�}_���J�5����g���r��3����d�#Z^��oM�A娽�A4>:�kZ46H�ڔ�ʤ�A���㌠��f�rs�i�1Օ�^7��'UI�ڄ���:������gWR���捖��~>��ێ嘎+&��3�nX�In��K���Yz���猠G�'���Y|>%_7�+G%�?�C8��$��>��hj�*.�T����j�J�/ϒ58���(�Wн���U�z�(��*��~���(;s��<:r�"%OjgZ���.�Z��39��J�תB-����k�oG_ �/SiY.h�"��͔�`�r�p2�zL������]N9|Zݡ8�ß�^� �0�J�\�~D�^�H�k7�������_��粟o:�W�=��]��8��������;Ѻ�B���F��:3-�+8	r�K�ǈVW�Y�L4�I���"���t ��|�VKu�74�ZG���EL/��
w8��|/TE�2�T��W��=��^��S �O�y^v+%�m��&r8D�m:u�e���>�%�r�-�O�hV=�/�/� �wH��xB8o����Q�?l˗�E_Z=�U"�A�ل'��<ƍR�>��D���m)"K�9���#)�Hu8R�6��Ց��#eI��f�>�!t#���'z7��Yj7k����d�J �CK�}|U�p&I��&� U^�@Q��JHy$-B!�Ҵ����Ս��E�)���@�!�+*��c]]]����[� ���k]X�eb�Z���T�s��$w����}�k����}�{��'T�ĪI��F��� ���5����?��ބ�>�U;\��e�����g��8����\ck��!��7x���5U9�ˑv��5\�%�#$��D뤯����Y�#�������Ғ�S�7`�1���Q��.�QX7�����P�,��G���~*��� �} m4������<��EQWh)w^���J7�S�����;�R�*�9VJQ���A5��*�O�!R�j�`�����-
{H{��7�4��c���@��%�/�����d��/�R��4��Ua�AXq>���!3Z����Z��hu2���X��}���:>jV뼾w�gb�9����%<
���q���-Q���- ��gȓy?r����7�-��njm��?G%�j��ߊ�f�3��j�S.�[y���#��^��r�5�>:[��3�X	�E�xZ%�S��B�OJ��Os�1�uU��	Ŕ������Sʹ�����Z��Yj?b"��ä�����I�:@S��j����t�L-4���)�|���c%�1�$6��[�j'������w���.T��a�F���zz��m��sh����O��\H��u2|��JWz��CD�o��zp>>�����\�P��?�7`L_�Jo����u�we�UQ/�v�y�����_sL}oe�&*��V��`PmV`F��?C��H�˅���I0>��y�~��J�ֻKy��"4���;��9�߃B^�A~q� ��NV#1����3�K�W1�nBƧ��Y�����ЄT�cd���zc
�Xܸ҆�i�Ҿ�7�������n�xe��-%n妯9�򡨖�=���߳�,�{�R��ļ����o��`ǌ����J�!E�U��+˧IK�sw�]��~�zu˿�������k��~:��ҫ� ÿ9f�[;��E���L�a$l#��i�@���Oއ�����8CN_������qGx�w��._�]