<��'��JjW�i�I���21�ʼ��{�w��u�lAQr��p0+S/��.���ȁ5��^�K���H�|GRA1g��F������j��2�옽�e-��9��W��w:y:�Ɣ��A�Ö�7f�6���q~��ht7����'����ǋ�)?i�t��uFP(YK�.���v-��������U ���.�Ԧ�X������2�ښ�],l�����}{���8���Q�āq�
Έ����<�%k��>����-�}��8,�<�<I���Y��´in7"0\�nr 8��-�$U��{�Gm�����wF�3������[Y�w�EBhz@l~��n3�b4�������K���Ū�X��E����K^���E��>�&�T���].���Uo	w�3�]E*��F����񉭝�T�>fzI��mP�͓��c�/��(�%��5ފ�JY�q3&�����'O�mj������s�N��)![Iu�%�����.9�Z��m%�t�Et�C�͐CRJ��"���zQ�$�7|�����Y'�/pB{�?��=�s�J���Pf
�C;:e�14�%��Z��0�J_'jzLT~��*�`�t+\�Xl�N�0\�R��)�v���&bc�ђw���g��N�=8+l��)��L"<��}N��f�.���w�����s@���:�p>W�,��a��~2񓁟!�$&c7�V)s�/N�rG��;�4"Og�PmF_܆u��6�b�5
Nr9�i��
��� �8+F]3 @"N��!(�C`lti�/ߑd��MJGe�M?�>"۲F�X��q�#���E*��v��JeD�<�q�}j���Cm�u�"j,�|��9H��|��j'Ӟח�e��<b����
^+Õ
����TbCRo�zb�avt�nD]0h�I�M��eZ7ϙ�U��N_���Zg}
���ի�l��,gϘ �Z��m��$g���6�������~�%�b$7߹��z�6;��]�uI�nꢾj+Z>e�Vmu��.
��������E�7Y��eSh�}���A�F�p��(�j/���KHx����6 �J�6cx(O��\j������X�<vޭr�<g�ǆ�]aso�0�f0J�'U֌�4�?��fM���r��m������8�K��8��{=���y�FE��M���ˇ&���*��U��5.3�Y7�L�\��U�`��Y��.Vöx��hO��<��h�2z�K�ȋ�d�"�����\mr�W��lN��C�-�!S�՛�ۊl�o�,HU�R�9ˡ�j��r�Tg3�R�j'bo�ZTF�,�lf�7S���UW��)��h�r}���ƥMGd�c�^7�\�f�r���5��9&�R-�H�R��e3>+t	Ø�B8�݀�S�#���<+��^�hC�G?G؝�T�4��{�_k0X��U��mf�B�_������9��R�ˋ\��23�	�p�hy��%��6ۑx�j��R�;$��y���ǦK� ��^Tr{|$��5���J�I�G_�w��o���m�e�~ʳ:����AЖ'6��^Ʉ�O���7ٲA���z!�n����X3�ɍ��e5Ŀ�Klc,��nŠ������/��#K�b�KXg�̷����4�I*�y�EO�.M�պ�&Us���-�+;`؇�ݩ��ZY�s��ݲ����	5Tx�% ��#��w��/W��m�6�L��[Fn+���*�Taeg�I/�_R{(ז4�'/Q��J��dԌX��v< �Gfɢ|)븍���#���m�������C$��\������xN�⚻I$���ŀ�	�V킺�|3C�c���<���R�{Ƙ��,��-[G�rF��jGU���Ӹ��U#�j��-3�cv�C��d%�X�<�8������a@+C�A
����K*߻�2�dă�������l�OR�1����1��k���buD1q�"Evu�h׆Rc�	�e�&��(��bu�E�s�2c�����=�J^f5>��O���j׿��\nq>�L����vt�8g=Kwe;�n</��!lh���B��Y�/sk&�ׅ�g=r;�! ;#��B,��MM���&ީK�u���bsrXlU��H�Kq>0]~n��cjCJ���F�"u~�ka�u�ް(RY��)V+���b�N@@"�PJllX����b�>(V������>��z�@ၚ���p�F-?�����oy�3��/Q%-�\+`sXܯ��X�U���45�� IhHl���Ix�ԣ���*a1�Y/V�Hw���ij}A���Ɛ��C�m0ǜ����M�^4s�����'��l�%�KA�YtI�v��3���x�j���a:����M�t��>E�?��E��=�'��h��ߣ�
���]ˀ�9�����OY�[�n�Z�����%q&�Y�}��Hfx]�-�/>q�2�ە��tE(ʀ�|х.?���sX��6�,�U��A,\�Ki�7�B%���!������`}�w�ٖ������J�}�o%�柿�!�X�O�CzI����h᰾�������[����Z���%@�ߨ^e4����C�B�29u�,0V�+.�υ��P�,&z3ы{ec��6��d�;b�,=uX0A�����я����0%ҐB��c>�������V�}K��!os����=;u_vԻկr��)�C��x-�m� '�)���Ih�I�s�G�� �P�%Y��ťݱO�vYz�;�����U����,�9���H��ٵL�n����ϕ�s�����1�F���:��G��D+h���6����:|�h����z���P��C<��P��.��wwڪ8�/´�],�IŪ�A|�)�w��Y;�l=�G�ƪ��sy����}�}U1�R5 UԄ��Ҫ@C�lFhU=��-$Լ��֣����-%�U4��$�b(��vg��J�)��BDdy��Z�o�ђvzz��zۗ#�F�^x���I�8G/.���J)%AO�ğ��3p~�rG�i�]�v�����-;N�˥�3����_�����pO�g�N�.�o��C�4�X��g���n��L�*C5�u�z24�gػ�B+�Y�]��&ē{/����r��Z"ʢ%eV�ç�$>���jݗ�W�h��gX��(�fGA�-��"7��άs���O<�P�ˡ�w?,�C���GKΊo���rKկ�+�Ln6ȲcQ��˖��2�M��/���9?��/7�Ƚ�1��_�����i'�����6=���ү��}��=οo����U�(��ߒ��\���T0m�$6�����KKRl�E~)~���3��N�S�v��˘�Sw��qf�4��]zw���.m��(F]M��+�K5%�!ޥw�'v�������.)V������#��m�-������^hAu�VݻM�n׽;��z�h��s(����,�K�F���~6�1�'��xr��p��Q9����r�me�YjakGE}Ipp�HA��J�嬟a�e}Vk��󚮑�~�L��Y�d�HgmN?0,��I�J�J��2�y�<`����t���Z}O�-��G�cZ��$��@=e�4Թ�7��)�̝[�}Do���ch�M�@r�a���Z�B 1�9sT��n�?R/�7{ND��u8��s�~ޮ���+�~i<��V7�D޿��?�m��������횈���k�ۏ*ep%#-�d���=ڌ�iF�7����~�9y��Qm�DH�X��c#�>��L�ÖEz�r�F���-�}5:�<�'pd�Vy�D��������m�I\r��}�2�!��s[1[[a=��xfVOp%����vy�[�
����6#�K���9��s��}xB��N��*�q�G����-���v�
35��]��pB�#��r0�gf@F�R�rP��9i"�P��D�T�ޮ���i�
��� |��VBh���籖������l��-�����/]�?3�X13|y�o��f�"ݷ@��ź��{��&~\ư�����2K܅��@Y���>��1#F����_bs�"D O\P���`U�r��i�7��q�m�غ�.���9��\��������'r!ٳ��+"6atCA�&U	��	�m��&�і7k#:��٘�c�!b�<ʘO?Ξ�X�AH��Qq]���V"�ל�D�4s��M�ס��e������p�=)\�gr$���c��������o)E2�:XW�RL�[�q�\� >��5��9+z��LZ�S���2.�~wG���7k�����.�9* *�-�N�z:}�&����muܖf  ��H���b���-��~��n�"����肔��r��y-�!�^�^���F$%6���3���L�
D��ܵ�x32Z���*�\�����f�͖QBIb����9�I�OxR8����&	�����FW����
�� �K]F�;|�˦�+LQS��ٱ��v���6e����5��*%����UV"�}�-���Yj��� 6���7�`Y��Q���eR��x�W
ɜ�|$%�S� ׮��Z��b�e#vt�;�u.*X>n�l56�U��4�h�Ҍ5���J�Y������������?s��04��_oe�!y�_�i[@�[I�,	H��զ� ߉(�@���X,�d��.yAK���Y=2��aYp�B�Ǘe�s��,d+W��fV���ci�TTT���ח�b��'��:�d)8�|��&��VF��6k��:�?�m"+��<oh)�`�l�X�1���Ȝ�%¹��h���,���W���k��s�dO��ɜ+�79��>W���E��v����O��4��h�ݗ+0�J�]�@��
̸R�YW*0�� ^�
��%��lB����AY��;x�s���`(�`�	(�g�� ��"�h�(��$��W��2��^�Owr�إ���0X�CM]"����cU��6]��G��S�i��'���$3_ot��U�#ѕ�.��]�JU�����X��_�����!���9m�{��>�%D�$��7��mz2$#bR��7&U��7���p��9��z����u�A��e��\!S��|��uq�M�8;���CÂ�t��gPn�qqނ+�[ˬ�m��~�nb�E�q�ʫ����woGΨ���Гr�?�r@�&5�J]hיYw�8��wx!��7�SW�`���! ,��_��ز���s���lj�$��������ϵI���L�b#~�k�)��m�y�ɟ�n�5�<:�+Lb�
�*��X$Y���D�h�'�ˌ�rM-�&��r9^A����{�詟������)��e�\	({ �\��F� 2F[�$ ¸%l�E��(IG�b?F\B���z9����\�T�
�<����,B�lF��#���lb"�Xu�<{��(Ve�F��{*L�S�#D�u�j܎���M�t��S�f��V�S�S���Y�`�2�K .b�@�6�n����3�n@(�q�Y��.H~�Hx::撥��4��[�����ܑ��p�
��v�$��\q��hl��V��+�46(�u�\ژ�Un-˄r��T��e5�#��9����l��5�*YC��#�#��O�(sRT�{N���m	Bˡ��Q�:��PW�����*�o��l�C&\�6���I��a(O�JK9�ņ��R4>�Jwej�ɏd���a�9�.�z�M�b�����d6���}��4"��-3��d����� {Yb��P�C��\�4,�`�H���g@�t�\:(X4Rf�����!�!q��$��J�%p��6���1�B&s�
Ss��Ĩ =�ޱ�F-#� f�dN�R{�p�R9������x+���=ZlzN�1���Cח�$&v��'?$cˊ�K[Z�uk~c�nd�J�ױN�&I�LP#~'s/K�,O�ߟ�T)#!:��2�J�'!Ni��e�����i�M���+c�bt�sL�U)Ѯ�Y�,q�kɶ�:X`i�$)�F�Bf��BL��I�:@o�G
��'��C����V�-m���2�I ͩ�x�@��W�A  u0X�����&��c��1H޿����� @�,��_ڶ%s��d�m�-5�`���A��f��,��]̉R�k73�)(�Hach殈s{�I�'�m�z�V��JH�m�M���ˀ}�*��G�``k/v�U�-�ˁ�s`{�