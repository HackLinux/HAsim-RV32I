                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                RIFF@7  WAVEfmt      +  +    data�6  yy{~~�����������������������������{{������������������������������������~~�����~~{~��������������������������������������������������{{{{~~~���������~~���������{~�����������������������������������������~~~~{{{~������������������������������������������������~~~~����������������������������������{yyyy{{{{yyvqvy~������ǿ��v^YYVS^icN9333AYs������ʺ��iY^iv������vNFYv���ǲ�{i^VQQQQ[q������aAAc����ǥ�iacq~��������{n^QNYs�����y^QS^q���������y~��~�������qiqvy������{v{ykiqsv����vqqffqyy��������������������{yy�������~{qkiifnv��������������������{{{{{~����~{ysvy{��{������yy����������y��{vy�����{yvvv~��������~qqy��yy����y~������������{iYQQQ^qi^YYQKYq��������YCS{������YKiK9�����S!#n�����݀!!!!!c����ݥ�{6.c�����şs.!^�����Ϣf6!!1^������ϯ�V6)3Y�����ǚvYKA11>a������vYA1.1Ii����ª�q[IFYs�����ŧ�nQ6.9Yv�������iF36F^{��������cVQYv��������qaYY[q�������{qc^^cq~������yica^iy��������siiiq{�������vaKIQYi{�������q^aqy���������vqvyy��������vYYYV[^n������c[Yqnq��������y�������Ϳ���ycQAFQ[iqnkcSQY[fv���~yiYFy�����i�����Yi������҅9F�����ߗ)!Fi������ߝ!V�����ݝ^1!!s�����ߗ^>)!!I������ϭ{C!!1i���߿�c6!!!!9Y�����ݟc9!&;c�����ϧ�[6#!!+Ca{�����sS9!!9Yv����ҿ��fYQYi����Ǻ���{cKAAIYv������v^A9AVs���ǧ���iYY^iq��������kia^is{��~{�v^SIIQQYf���������{������������{���{��qIKKKY^Y^iikkccy����Ǣ�������ǗYv�v�������K9S!!��yF!i��~���ߟ�f3���f�ݧ3Y���V)Vy;!A��vA�͊IY���v�������ͧ����v��������kv��[ACQQI[qvqnnnqiciv~�������������~y���vy�qcacii^Yacafqqvicckqy�����������������{v~������qiii{���{iYQQi��y�vfk��������{��������v{������q^f^I9AAIckYCKYaa~����������ǵ���yn�Ϳ�yyQ9Yvs{�yinQ3S���������������c��yv�qs�qQcqaSiYQ{�����i)!!����߯q!!c��3!����i!!v����ϏI�����ߏ!!�����{!a��s�ݪY{��{vc��;���߭���QA~��s��ǲ�kiv!!Iy����iKQKA99Qy����Ϳ���������������iK)!&A^a���iQA9;1Qfy��������ů���������sK!!!!!!AYiviivvcns�������¿����������vciYAAKY^[^cfy�vv��y~���������������vqcQiyaIak^c�ia������������SQIFAcQAQqiy��i������������!C9#C!!!V��������寏���⿊��9!)A+.Q�߭y��������ק�ק����qQF9!!KA!;9Y{������������ҷ����vn^QC;A;..)!!!.AYq�����������׿���cKY��y��ki[IS[^YNA3+9QSYy���������߿��������YKI.!&)1FYYqyy������������ŭ����~~qYINFYFK[QQq^Y{�����������ů��Yqqa[n���qnYy�{{���~�n[ikYKYivvYQQA.!A�����n��y���F���13�������v�����	!i>Cq����������ꀲ��ݿϧ!	^Qi9I!����ߧ��������ߏiKQK63!>ys)!;Qi������������߭a&!��׏�a!1a��{A!!!>��ů�q9!N�����׵�v����f+!!!I3!!9~�����������ڵ�q^YKA>!!Fsvqiv������Ǫª�����iA3[����ǷvFIQI991Iq^CAICi����������ҒcQ9!.!!!���������������S!!�ǿ��