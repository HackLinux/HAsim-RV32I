�f�3��PV�澽Z#�T��f<��ƚ붝}5�+{�W]��]�e/�uX-%�4�hMj�ԣ�|�q����b*+�<ge7��u攉\^�M���l�c����������L��%��[��1Xo��V���e �fb�\a!rc���r� ¦s���^\����7b����[��F�D����0���h�[���h�h'��xw'YǺ�\~{]�*�d��j9!1��ē#9�MQm�����8����4��[���� i���de���U5��lܑ�I��exd��&�@��P����ҕ�RV�����ܛ(b�VӅEF��e_�{X�2�N�cf�U?h'�IK�Ǧ�h����`���q�(����Ժ���&{��ʍ^~.s�k`��p�wK��"z��K�E46~��~�ej�۩�����h㏀�Rm�Ad����xP`�.}w�y�ͻ�i��/��)}�c_|��O�⃷  �9��*��`����U.�DW���T���qV����0z<Mӌ!�JR�3^`TbZ����'��}#�(I���U�9�{ܳ����Lf��Z"<�pU�&��;K���s�y��,�Y���?8�ҝ�d�4��P�QH�m�<�Mk�W��G�.L�A�s���աp�n��qē������a�C��9=_Ut�Suո���QW��|��2U4JǰQ>��"4�L�.�q��[~��.�A[Պ?���p����M�u!�n(Y�t�����E��|�H�
ލk}?�o����e*��㚌&�{Ԯp �2����Ldzn�#��`Z���AiF/�'��w-�~����������CߔiR�0��6S��O0��{4/�v�Ӽ��FRQ��|�jK6֡SA%�⹂A�a
NN?eaǒ��ѷ��+�w�e�fD��G�-�6�U���(��å�PZ�
?�������?�<$J�{kD�bd�;�*Xc�
lSl"�������	�v��zɚ2:!�æO/"������e��@�[ui�	T��(74�#G	Õ^����(��k��a ��wf��ؔ�]���7 7�TM�g�#�Rgt\
t��9�rm[+My���m���k�vѫܯx��c��D)*SH*Sԗ;򂛴��³�Y�4���s�#�F�>�	�ku1TS�Z���"��ən���&����U7A�1���B[��)�2�j%��S���!s�|�T�_;�N���J���Yab}�v��OC����k=>	��xx�1�"���fkک�E�X��1����'f�����ԎZՑ|c�s�V�$�M���q�ؤ�3b ��bx�	T ����/�8!�%��~�4���k�cHբ�f�z������m�G���($�H�d�Sad���a�X���`>��	Ј�$G��(�Eݖc�m6�'����1%�-�+�1cP��1��fy
��m�Oi�,%��Jܣ\�_� o;`FgN9F!v��=w�Ej�e&�-�OJ�^�[��Z
����I/�C���]i���w�C7]{����v�l|CRL�wuؒ�c��Ő�xe�ϫ�x]���G@ᥭ(�]l��\���*�%p>+x;1X�կ��KTE\�K���8��7�4�tr�������^"��8�5�~�z����B��FTʠ��J'�)�b=�ɚ�b�B�Hɔ���*���W�&ߠ�q�@�A�����]�y�#�[Q�,&[~0{�	r�ފ������w�
4O�4�"�"�4������î�hi��7�k��s�>���6ɷ=2LL,Q�1������"L�Ӵq�y��>nK��_K�� l��C����k]��"�;G�u7�)�_�h#ј���ҟ�O�hOJ�,D�*%0��X�o���هvj[I��}%qc����N�*F����ӷ���h'��B�ҢN�pe7�O��n��gP�ѳj�l�=9p̥����t��L;/���e]o~�.��RwQb]�`�9يV%Ǿ�˜y�"J���D����;M�\��6���Q��T6�Z���9�+��E��y���z)��(�����/G.�v#i�bp4ܐ10��m9�ڮ��6Ѫ�]"ّU��6Q����4�\پ)��z�pek�N�v�;ѣa�:;h�hk�<��8Tg�F�~��~�@%���9����o{�*�&������dTo�.B�Amȡ�s�f�������y6az��CzY9*�����z����ݸo[W��2�Ec2<i�h};Β?��"Ht��2l�J��$f����0t��>*R�V�OY��b�݇��@!U�s����	&f��c���[T�+Z�wmVg�" �/���B���P��W慨���H_3[�1Ml�}� �=�J�Pߑ��y�DpAzx��`p�
#[�:'��tޖ�b��Vu�݁) �۔�~�1}�͗&�����) ����I���!�w�?  Pe��X5�Q�[1��O�2�p%xAA�^4�ޯX��g�G�$���������P >�OK���cp*�!8��i�>��ސ�T�4�jɏ��W#��9���d���,��#�}N8�܍:y�%ڹl�5��-O��	? � r�@|=x����*�8w�H��[#"� ��N��X�[���(��`Z�1t/����l��5���2�R�B_f��by26˦�@�>	����Q��a���á��<ʹ��2u�9�<=��	�	?�KQ0�
ڷ��C<�T7@p� mڃ�_ʵ����;��D��֔Bl?_탔\��b,ŏ[�)c�>��k�jf�m����3��}5:P���ֱ���Sg���/K��(�ﱦf��~���20��l�ۚ[j/�H�aA�M��Ɍ��;wg;7��"<��U�^i<*�A
3�P��wTK'��ء� �D��5GT��h�b;�1�79��N$�IrމY�2�����h[O��w@6d��6\]�,���l�Д]C� ]s|���l۶m۶m۶m۶m�v�?�&�$���[=�S]���,g�*N���_�_N^�"LDK@���f��h��JY��7Im�-,�eo�B�v����p�y|�Я����b|�rc>�� t�KK���∿�RX�����6r���_î�әQ3�2���E��?��{6��<�!/��{D���p&��(&n�a�^�aC�C\�P�8v���	���#D��G43�p�`�����aD����sE��6O,�`�h���_���L�^���#@{���KG�>��/��4�����3e{c�rB�6��ǭ&�Y��ʟ��ӊ�#cL"w`�1Y��5��O�5�ԇ����Mr��r���'rɰ|
���p�r�ox�;G�0�~	q�א�ȿ�B�_���^��F94�^�|�g��~wRϏ{B�d�B�Y{[�/ x�� [��^�^���r�T�d��/��r�yˤ}N��}���|����"%zYY[��n�\_up�7d�ym��#��WqG�G���7�$O�VEWL��~x�@86���D=��Po�T>{8+�a�[�ѵVoRU^�A�I��6 �p	!!'�%tF��B��r���RB}��8�D���f�m�wV���w����ߞh�x����v�?D��r��P�v|�r��h��
1͝�o�ԒIߠ�W[��������%f�m�f�*jT��Q'��h���>/���͸����Cp4Lh���t_���^�"@&.����4)ş�2]�
z{�����h���miis�fo��Я�P�,�AC렶��EͣGT�_��t$�2��,;��`�޲�2��]����XY��g�:�}���yr���b���jM�'��}7�g�F�"�?D*��6)7�	�b�`�+ZJ}"Z޵�P�vnZG Gkl:F���w�]��U�\��O(��ù_����=@��C�����!.Z&\��?�������)�?^y�#�,��3�f���M�j/�30�#9]Y�iA��
�?���Dܿ�`A1����H��#ܕ���(��S*׽����ջuu��Q�.��5��������I��~V�!r�E'K�0�!�+fϿ:Y�gs5����x��S��^��&e��J�#$>ΛB����r�w.?Q�~�������#VlMh�3�:���z�f�Ƅ��ލ�hI-���}��`Ԛ�4G}T&����D���w��9�-lN"�����Yv�ڸj��m�ҡ=���Pl�<sR���IE���	�S��c��R�	�,�S�R�f���O$�_&����"N�H�	�ʥ��m��2v���)~���M*8���0<%��Z�H�f�O>���|n2b� ������j�����sk*�~ �-8K%��;���-!�B@�_z���5=q���k/�G�Ϗ��������pA���M�w�y��"���ki�;	��"=K��m�#��S8oy.��+bE�?vb��D�����oG�>h&��Id�z�.����,���kX��(3C�WS��brnΈ�Z�-R�����;/��T��kIv�m�s�>�{*>f�l�ӷ�p\�*H1�i�N����%g�zH�����ۊ&���2�F�M�
X�d��XƟ-#�=(�-8�F�/���CL�Wcb��x#��u��8��N!S���0?&tRR����I"K�ٲ�S�"Dh~<4�-����8�����aj�k����c/M�Nx��'�w��$�p�5�O�Wc�9�^��ޛh3V���>�Xh�	����Ta�Ii�
�8��.e��y�Z��-��b�S���p�΀�y��K�B͡�ȡ�0������*��],mFYa���v\C6���WݮG'�]-_w2����	�����3^����'����>�βc��?5GN�����/�c7��b2GN��i��I�\r/�����4���W�W�adN�p�M��a�1�1�`�n!}h���9p�䎝A����e���@�W����'A*�����n�W�vS��o�g��].۬��l2w��h�7a��ʓ�c�_N��w{< .�S��~}sI?�X�'|�W� M�[(�>�}k��X�"Ef�q.������p�����ȬE�Z�i�ħ�������������=G񏳂W|��`/��8�1�&�9�*�K��P��]AT�� M�e��|ڡ�x��Ӛ�i�8��g�$8��E'	�oUIM?����,�&�8_�"ΐE�&@QQn����Yz"��@�V�F�KZy�9Ȉ��U���3`5+�Q9����xÌ+b����v����}5ȪT>:�~L�<B���r(]�쁗Faj�:0r8��� |�G���l�D��}l&X���<��7��ͤ�?U`*��Zԓ�{�����v�ǩ���-�e�?��H��aޗ"Hש����D��[�t����擣�Nk�ʦ��K�b�@���.�">��.-�ŝJN���ѐL��o��Ӏ��-|>���*C�_��;�q)�d���Ҙa�+_S:��J�XĽm�4X�;%�d�/�R��!KS������ɻŗZ�z���[g����� ���Ӑ�Y���s�X��o�(u�>I��]����P&�w�߱L�(�6�j;��6��{H�A�>e�e��=Xf�S:��V�-!D�ۢm�ꑃ�����-M�����b��O~�"���:��L&�G^ɓ�tf�W��va���g��_�c��n$Q��$gplu������~<��^�|p��v�3��ߔ�;Bl\�cbr7��G�5��C춤�/��<_Y���bw�����e?�B����u�T�p\��Dͩ�]R���;`��ԑ���Q��{�h�Ӊ�`΄Y��Y�*0��{���i�I6���α[�>4S�T'G��Ax��B>���摊`��ճfބa�^J/��A��¿>#��p���˷S53e�4<.��R;i�C��r����-�"�Σ��棷��L������*��'2^�UV���C�Z�����{��?�N���/P�b�����z*�=���'ɑ���}c�=�0n���#���x�T6�n�}�����u>9�o飘i�p�c��p�0m��f�K�Ś�V��\^��Fޞm�j�&��<�Ȉ�@��������4�+@b�61E���q�[��?�V��m��N��L��	EI�&�lsy+v#@�ge;Y�6���i��i~��Ady�>�[P���G\Bjn0T)�u�$�3�2�eт84�Z��a@=�'�_|��;ϟ�C�|��ݢY٤����mi���U�Ε�̩�
r/V��W7q��p�K��SG�;=�&��Z�/?�����v� ��H6gʓ�@2�,NR��ayWt�=��'��:�c*��$��t�W���	�6�-��y;���«���`���t��&W;�P�{]N�K� �\�3}ƫZB2E+���s��4Ü7{�r9g�9߰�ϱrh-F�PZ�Ȏ&��j�ց���nPUB]�Y�@�T'�z��#T���� ���=.��kB��3�oJ���܆`�v���i?/ب�Ȭ�-�}Q��&�r�'8����#��VF9�,|p��?�.��=��������H��u	َ\D�ױ3P\��z-���Uu@J�<�c�W�iz�{`�z0!���d;~G�_;�l�R:�Ml���a�s��~j+$ܷ���w$H�k��k%����|{�M����|�$%sʺY��`���L<�e�g�A��b��:������Z��zaE�������:�Rb��L��O���
��Y��1�H}��F��Mޡ��Ҿ�k�l�F��HY���K�p���߻'�S�z=�8�P!2! �!cC�q�!�X��@�Pj����� 2�e4��$�֤U�)>7<�qJ����7�_!{�a=���=�c��9�9�t��j�{����$2�h?4G��k���-�K��n$F$y#1��`��V�FW��(�ǜx�sC�l`% B�@9�>V�j�,�����ɷ�(���{H졀`�ڎF�=%�uv�F~�/U$3F>�0�����IYؙ�]Bz�Ǣ�cE��.	Zq\�P�ŭ34_�ĲnĤ9��{]|�6��+>�Q�P�&�L�N����V_��2wW(7��q���&Ĩ�C�@G�'�R:�{��؞j�,�wY�S;�B)sS[<р���r���.��:x�K�v�*�;�G�>ro��=rP��}(�S(�����GL�jOQtc|��o�tm~ �z��"�[�L���'��m�?u%z�_R}0` p ��w3�w�p�W��,o��}�n '>%|+����}�wV�_e�_�`�R}�R֞��t��x��JѯŅ�O�p���N��>s�;M����=~�m�I��%^`���ןN���X�G�ߕG	p�r?Ou�,�BY����o?�BF��w��	�љ�G0�m��U ���P��ݗ�ĜS'~�|W�y.�s�f9�M��}���d?�>���v�w)T�WSr�*����ڏ-v�h�]~�ZP�BءR"h�&ͬO$�zHep~�Կ@�hKG����X1V���S�2Z8�9��XJ۰�����/��b�b&:;�S�����M8z&���H�E�ӫ��W�<�g����3Ur5�?<��� 9��7�T���򔃃���i��؂�I9A˜�F'����S�5t�z��W��c��$�s �E.V�#\�q�9��t�h�U�co�i.L�Lo~rB)��b����ar<�V��$���%7!R;.�n���2(A��>V��Yi��������;(1�J��<�9��A�Ww;�b&�-8/����H���`�<�]w�q����n������d4��mI�d���T^���� Z+.�K�&�1�+\0̗���1��
e�U�M
AӺ#"�����Ue�b�EС�p+:���{��,~T����qSpǈG�S��
FB��m�I�!EK�`��W9`�5�sv�{aW0��½��ʔ� *���i�`�-���j���_�e_k{��(-��^��Iֹ�XU�6$�ೌn��х9�-�٢�p�A���@�d7f�;��)٘����mq?��9i˹��r!��԰,��k_m�C���IP�L*.8����댏a�撶
�]1v�� �%-w�A��N�[�AaUr��:�^���m_۱�+'3�۔�hw��#�j�ߕi(���ZlkG6���&����Χ����B'R���ރ5���Be����vTC*W���L&5�l㖸�T������Q�z9_����HssKB|���amQ����g��մ� �=��V܂Q�44�<R3�������2ՋŨi���?�=��
�+ޕl��L�.a/,��pO�8�I��a��WГ�3s��8УG��BC�df�W侂�O�d�x��OV�:�m��G�6�mTm17��7wf�6#�<�ӻ2��ӨҦ}z�XSԇ��m��,�#D�H��`�"\���>����	XL���Y|���'�SI��|�?�+V.�6��;��7���lg��]�K8��Ě�����AL��&���F��c�Ic��M����$��5t�^����7�����i2�{��)T�mp8�m�dPS��9�)�O%���A� %X���qi�Ic���`�MӍ�u�4�aV��#4��q��#p���2�ۺf��I[R�gV)<�+�֍��T7����:��{���.X����I*�f����մW�J,�غM y��I)*I����pb��kg	���-K���	�`��%�[���_��$_�MIkDM��רI D9P1���ӮU�� %�x��90�~�KZ��|�M��n	�l���^��{�{��-��<;H`�I灬U�t�ې&==�4 c�çS��"}z�����kn"0Ѻ��SSNG�y'�!�h4嬹uE��8�U�����-���Y�&I�'+�s"�t�{�ʒ�I�����j�C��(�?eXc�KqE]�f�����q�Ѧ���f�ܬ�G$�-���,�wq���Ν٪P�M�PgE�Sl�WQ�X����k�5�	�'vbb3��ܳf�!���x�ѩ�s�-�S�i׏H^2�<�ߖ�\�Ű�G��bF��g�_E0k&���e2;��>u�T8�(4��`Fd���زx�v@����Ã
9Lp��E�}YS�T�:�\ĉ���D���R$���i����Y����Sΐ�aUDɨs��}0��G����.d���V8�`d3.��S<�%&,H�~�>;��狼a��/rɯ��UZ�!O@<��8�-)R�E�\�+�^<6�6T��N�`U�l���A�i){��7�s4g��Pa�����;>bX�Ap��h��V��޳W��VpK����@_R�[��ޫ@Faq7-C]����;�=��E�q�?ͺ����o�m����6��h�F,+ۺ.x�*s��j�����g�������M����o(4�oO�OP/���:��\�����0�"0��M�k�+�Р���ːVAym��?/~9k�Z9+gLr%�=*��Q��gB-�7ΌF@|��Bw��n|���͡��Єzۻ^�ժ�z�g�� �:~e-��z�H�%X��6K��XԇfO _O�(s2�hh�eA1{BO2悪�,gfW��m�3u�8v�Q#��cǻe�^�L�ݖ#����'F�s���(��v�1	���Aj�W,,��v۝A6��bV�s"g�^c���;E,I�8T��!�Ί���T#}�7��o�'���Tb�1��E\t��y*�_��+���s�^3�f�[���*	
8�j3'��@Y�pV��v}3J��b����F���'Lh���"�"m�K޷M���q�n}N�?��yx~܈SU�0}�"�\�h���P�@tf"�Md����E���j���z��\��ߦ���	[��%E�T|�٨={��{3-3M���%[�O(Sj�ɝ�nW4�����%4L�z���݄�0���bl�K��T�����M(�i����Y�KZ�4��C�F�tM���ʄ_F�s�"�S�GK2�jR��u���[��N$y�j*����%�&�|~wh/��%�O+�h��ByRqi[5�b��G]�hz[N���b�����
�Ʉg�4�c���n՜d�:5������#y����~�|���#�Ln
6G�bl�'a)��T��6���3��Fg�<�5S�c�����ZQ��W�h�l�G35����v�m�˨�J�[M���elϜ	�e���6������ޮOsY�6T%'%�-����vP�-K[��{ԋ�	?^!�Y��L"��1%'�M!�E��>R�������Ϭ�Vw_R�>�Z(8�J���Y�v6�7	��}���K��
�ێ�C�F���hG�3+Ox��<�;w���~B��ٝ�'��嬛�dj��5��M�����.O�c������\��F�"6cd���q~PW���-�Ύ~�ο�%�;��;@����3�W�  

����5��  �螝��'�-�=����6�0M҅:ih���Yg�n������<�ӂ�R�]L1�X˚��Ob����p�	-�i��H�Ɇ�l����)��6;M��M��;}s�s���������Z@�4�sC��۷q��ĺ�N����R��OwJ��z��ܺ.���O�P&!�a���|��Ku'�}7kr�I�����x`�@h��K�Sov�z�;4����?`�ꛇEy�q'`�i�A�s�0&q�,����I��j~�q��Gb^1>�~7�;]nnK�Z�~�L�N�lY�J ����o��X¨��2��<��<��?p!��:	G��N�Ĉ��B��3�ə�ۇ�S�[ϴ��c�2�ϭU2����l��$a`�}^�gԺ��LZ�+Ӧ_pv2��;Y�O�zv���jӯR����D*X�I�����W:�Њ�b�-��|���0SEH2�b��r��P�]
�R�z,(���yV��ֶ@Y�^�N��>A1�����D/7�Ƞ���E�Pe�^z��}����..����Gm@� ���;m�t�C��^s=w^{<W5I-��j+���*3��-�j~
6s��ڦ!��x��.)�;XC,��R#�e&0�>6���uF�@0�vn�	�㗭���`�ô�7�܈?��L���i#��gg̈́lN,�hbnk�c'cA��qv�,Yp��`j̢��'��.���X���쩶T�ǧ�'��B��`�m21(�V�.�)$���9��*Ow<�2�'%�kn� ��~=3��ꗠU�8�m�d^ �3�y�Ri�J'χ
*˺C�蚌�����Tރ�~��^���F�b3Vd��Dd)��N�v�����\�ZӴ"�h����0�\mE�#ikh��S�Yn�a65�f�[`�����0Y�G���֊j$�&+
S�D��>���p�}���}N�E�~���#:%}?Y�eAS��]Q6��~]�8�����:�:���p]މ(~�J`�u�~;;5�Ur1:�Ͻ�do��Nb������j}p� "X|W��S,p�37�%�`��6:�~��[��lwm�xlϏ9��?Ӆ]�<c���y���;*�lǳĶ�W��pҫUl�i����Rskc��=���3��  ��|�Wt���N!��d,�ź� �=- �ۋ@��G�0�CY)��yr���۱]��6��e�����8�ؘ������gG��͗�������'C������`�
�ti�񄒓�/ �H���Յ�����<�(+!�ViP����U�`�P�Bpc�hVS$8��9�E�/X�6���cL�_u����޳ԅ��uV���Aj�Yx�����Oiu�3�q�\#6�)Y_�%]4FW�,Lή��6���犵��"a)wG��d&"�
�5_j(>��1֦M>=����7��2��}TkQH�<>24٘VP�&Gq��c�y�&	_�pS%��Y��ٹ�S�z_�l�оM����8��پ���OdFf�����#D%���	��Y�%��H"�D�ϸPP������j��)!�(;J�%ɋ�p(�kB$ ���Ѻ$8�ex�)fǟ���a��O�޷���Ե�Y������K��3M��E�IräV�rD<!�HԇͰ���iC��旎yefIEd�.���	�0,J/�����(.'L��J.�ں�ZF��;Տ߂����jVL�z\�D�r6�mb�	|�]a�V��H��&5X:�V��)�ے����Z�����bC��ѻ}Z ��#��M��}Hm>�Yt���{m��� �c/�i�Y� W�h�����U}�a��.���u� �GjT�xOy�oh��}�����6 ����L��N�z�[X�!��tψ�Х �!?�t�9a�>N�;h�׾�h}����z5 ��W%D�����~-@u&~7z�h���?��_h� �7�����>�h�`��t�x�J�}���U(�3��g�����Êc�e��ÿ/�r?G�|o_.9�t� �����]5@��ׯ|����y�	�2�\M��78�e��.��?~�+��_-
��
�?w=�J��d��qw�xV�W����E�ߤ{=�EA�?9 ^5 E>@eB/�a·�߿b�_GE0�=2��9K8�����*"O��=�ϯ� z�p�O/D�			II	�����s-y�١TгSUS�zn��W�@�u���`^�B�W4H�*nE��$>���n����r���n�N���(k <�>H���ʨ\���@��.��F��� �_����{��hn[N��I�<���
��!w�(ţp�����d�V���,&���J�;D֕�HU�A��r�ۧ���f�5Y��2;�λؐ,�8^�M�w��0ۻ�ҙ�ٌD{+=O&��2[B�����A���9=� �/�,�)�L��$l��4d��� ���$e3��'�����ԙ�*5���Q�.�w�U���˳,;���G��!�K=D����&76�2I	<Nd��?m£X<���m�{�&
�鸢�v�f��n����Z�id�1]��0���,)�d�4l�Si��{h�[^aP��a�)kz����ς{���*Z|fʜ/��-ar�)��w����!al��b�܋W@��lB;T�У��@� �5*�S�O�6���~�U�.�����CS�J:,B�D8���->���I�`�s޴�%���5*�]���]h��}�Wx�)$�T[/'�ƲnB˽��t˶#H.��*+.���x��'hs
 yn-�	��s�[��idT��D	H��*��m�'�8>����%XÍq��L���/BWI��X���'�9pfCo�$���X�!�gy�H�X܋�㴃�$h�'���.3{�x�+����*�Y���)�K�> M�e��x�0snl�,���A^�ޗ��\�b' fSYTÂ�@)��
vD�;0������`n���y2�l<ji9Z�@�)�]���'��K�| ���i�?��Z��(um^S�FzЧ����[^��9�������������'�o� G���GU;;d�a��Յh[�x�5�Þ�Q���?���x��l�$���0O�I��wC�\�y���0�a��ho���JG�i�9xdh�L���-�oi�9��9�=�ΆP�L��KC�fb��7�o��"Qj�ˢ�	<�b���|��k�)B�7V��rtR��Ee��S�D�H[�ЅC����c����Юg�y��d�bn����֊��R�ڇd�oLF�t�Q�F�X�=��`�[씆�4ج����l*��Y<���jFY��+O�4�b�.���HzP�+����r�$O�� 9]t��ci%�G��Oe�++U��=��x�8�qiF�ul��Dic2��`zʼ�=���c�lE�`��>��O�8M�>&�V��:�qe_k ����*��I�x��#f���˰���� eґc���~��)H���Y7&���7z�rՠ�,�i)��E���j|�p)*���ǣ^<��c*e@X���Km"�d��?�mAn�z^s�;5���d%Ԏ��H��"^fR��˅��O?�`"U �0��O�d g��k�i�i�X��GX��,�H>X(I�B�*���$(@/,�-��?G�RS�"���'�Əf}=���;|�[�d����[���τiЅ�Gs��<�s�߾ �鏚�"�?�C/��+F��� x�.6QY�+!M��(���$7�3m$g���b�r%��:ٱ0!
i�g=q�Y\t�O���m�2w3S\
�ށ�����4Z���ϔ�3pi
�N{���hfv������-��ND����^��'�TSч_J�r&�5_�w"�)9����~��J�)����9�6@�Ga�M��T�ۛ�ȱ�I��$d�~�6��F����O�p����z����i��Ʀ�ح�'f�&���R��?m��V³�Z9r�Na�'D�l�	"2��O���]�5.�G�W�/<4��4��*&+@��ܗyĈX��r�k��Z�ٶC�>���1��g�u�
��ƪOG|�L�����q�Da�-� ��wS�Ӄ�<��B�z>k���Q ϝ��"��yw��\U#��k�t�'Ɗ�̂O�P��b����q�]xAi�t��.��0E>�֊�Aa*-�C1���b?o	�[M�YП�5 ����jt0���実�) sKr��7;�j��҅��AE��G�E�o6��w-�N�Qf���o=*4`J��B*b��X~�l��v����Ql�)-T�ep?���~g��QX����cM�F�C�b�'�>�P=Ք�F���"���h/Ϙ�N���2H���v
~�`�	4���8�mN�A�P)o�p)���#��nP0xK�0te'VC�,�y�^��}ܘ*܍
.X������a�vR/�ZC)2Aת����P!��5vc3:{����q!(�^���\�e'�	��H>J � �Z�ރ�G�d[E.���c�^�pY�����MȾ���0ʻ��EX�q��p���^Q��L�pe����v�*��z�r�bdG���Ҧ���|�K��c����U�U@��`��Uc��*�穬`�9�ִ���W��xCQJ}Ҝq�ª��EL��maL��Ci�7�
�s@ĪN�hYƣ>ː����r�����k]�򼻥���h����`�����s� g�46�l��.5��oq�t�y�����}��Y�\
g=Т��Lg��,���'���Z��9�\�o�+� �-�"�b���Hy�Y'��\}���N�A,�������g?�y}W��/2b�~�D3�jWu�7ʃ���	�4%X����RB=�R~n��,r�#7ɴwk0.U~1��	�;-�U����*��|�Lceu-(��h��M	�1��d�,͜3� �~���G�|n�� �}�&�᝗��41�XGfK�O=	FM�A��gt�� �|�����2UDWu�Բ��@����-s����6t���S�����KV7�C}I>ER�;%V7H��ؿ%��Iv	����鿷�߷��Euo4K0�F�#`������O5�7:�ǽ�%a��y6��Ka��M���nt�Ά�����M����-Z����P�ݳ?���������m��͕��w�V#�����A�����c�s~�{���ӧr�����6׳4�Ւ�����֕���H�m��[E��g��:�x�q���RE&Z�c5����y�$��6�[5�
 #� 
 ������fw��s�g�^�J�p���p���������7����˷�;�z�A���#���Dַ�jvҧ�ȷ�L���a�A�}�M�%����9S�}����<����W
�+���}G{v�����u�^����;���t��v���
���X�����b��������������7d�~�����w�}f|w����	���������|v����v�u��w��7z*�����OV�{c�o��q�@,  �e���6ݖ�P��ؐM�ExTq�#|�@���D�wޛ%Dl�3|��RVW+�o����N����`4�H��m<��Z\#�Vf�*��,�>��R��{�/-��ne���A�t(-�G��z�v�Ǽ�O��p4�^�~����6��Q8���g�k
^�Gy<�f$��;G��I��� ��E27���$z/�����&.�;�>��?�
_^���iɌq0��'�Z��Q�] +Eq4�9-���-�>�������� -@���H������
կ����
��#v�tǣ+O�e���x�<��:(Ⱥ-~�3�Xs�Q"�2����Ii���C�Da��)�8�i���<�����>i�M��R,���n�No��սC�$x�+S�sh������aCUv��%8L�
�i�6P�u�_!�ˀ&ݵ��D��	�N��n|?���uG�	��W_nZ���0���	Trޯf� �Z��@, ��\G��=0c�~��o�����nXx�����[ϴK9��#��J�ٿv��	��e}�����v;����>7���{aC���d����d�w�{�U������o�m�W	���K�F�}�o�/"�0�D�
��h����,k�_�[ܘ��ϖo52~�*n�n
_UBN��Cj�E#y#�
�$�U�8�k�n�N��~I�,=J����,�$n�c�S�Ḣ�tC��l>`��}1 k�i�}�֎��#���|�q�NE)}f���c���f�T�M��c��@eGkE�Z�Vܹ'�Y~\1cH��<ʤ���'҃��d��2�~z۠=�u�$L��qͦ��4��n�?�ղi��D(%���&�Y�j:�2�b��z#�q�S���>؂̞�WLz=��%�t̽=4�eN�0b>��%�vX�ՠ8WZ�^p}C��ƨҗqЧ]�\Ǚ op�A����:��ːI�����y~��}@*G��z{�@AT�����6M���(������?"~1�4gd�P$Ӯ�A���R{o�4�|�F?��{?�XtE��V��C��k��lo�(��'�#u��ı���O���h��#��g�ܜ�;�z;!��T'��:�~�b�.f[?��y�N�Aˑ�S�%T�cO�=$|�
I����;��ɢ�%R\]!��^� |U�?�g*�O�b�� kA�CD��6,+=G$)(<rA�"���S3��!�^���#-�)@t�>�6<7�"
�fU!D?���F�8)r�H�u:��I�yB,�$1$�LO�J�ky��P�u&����벪�<���-D���۳���*�U����#�%�^V�j^�=���{�b��kW�\�ƒᙕr���Z�'O��V2��awO�N��ZX-*���������Ta	�ouSZ�k��G��d=�p�g�d��3(ׇw�
����&y$��:����cQ8W�Sy�m�<}4{�8�������G���ɇ���?!��ɫ�D�B^I}+� � �X�r�as�tv�HRY���j�C��b�uTf�t9��8a*�,�[�r-�9�}��/�	�&f��̕`i\����uq2�
�À�A6x�.n`d�`�.��m;q��X��a������Ě���]F��?�٨B}zP��%��ی 	�T	�܁H�0��޶!�`Q��-8Q�#�V2�
qv��ʅ�a�nO�f��m�A��᪟��X�F�M�.[h��!���//��^۱�0��������N%`� �D.tV�p��[�^��&czm���U���uo2f��|Sk�����˘#��A���41�>t��<fy-��^f#��r�|/��
O`Z,_�k�E�B����T���E�"�Cg����fo\��uFZ��8�6�u�!����\��?��@�<��1���+-��� %�z��U6q�Ӝ����/䪦x'Ҽ7��7��X 
.aJ�^p�:ldx��
�k-�e'V�Y�Cj���4L>�|j�\�#���B�l��G�f��`�� q@]��hm�r�S�����F�3\~��؛Z�_�hml8L=}{�n��}�>����ӳC�Dؒ�X�������J����)9��D���� ��l���E�E�.J"�|��
�`��ӓP�gK;B�R'���$���{��ж	�C�*�Lh3*��Kh�oa�E3���Y2tW
kH�{�6���,��j�EMT:�%��@/�ҕ���6�^�@�jF�&�-�Psu�epn,[��v~���r�(%T>��$�l%��]�7���n�n��D,��r>�w�f4�����w.��UM�s���n8[�as��.'?�J���b�<rMB�($N8�?��o��f��4�s��<�F�,�J8��>~x��"��\�Ρ4��|wY*�uo5�0�oݑb �{�>f�q�+�-}��op9SFOR]q�ٷ��X� �RZ���H3SO�X�O9�]Ņc�e��M��s)�i�9���?=T�����Le����~�v��v'c�\mwm {m�}n��Z  �����u!�0q:L���j����9�ʽE,�P�U����f��a����CV(�!�jŉ&B����H��y"1���H��'��S��1���Fg�M+S�S��g�'�4!�j449��H�iWˀ���@�`eO��AY�W;���N D%�p�;#�&����Z�2>���?s���J9�dt3nLg6P	�#����(�7d
� �M�ףJ�)�g^����Q�L �R�ź�6��3�O��cL�n/���`��[Ś��G��8�!�:���8�YN�q�9��܄"�v���_+�$8J��c}��;�Z��y!C�+����T�+'��諵#�*�H�RѶ�s"�Y]����n���UW- �{�A]=f����GI5��j���<T�,޻�Q�\��M0Tzɇ�h�1�=��GO���� K�IA�=
��7\�U����&+ڂ���.f���v���:Kԙ��u�
�^9�+����K�!� .]����?bR��&?b�Oӊ�e.R[��?���Hq{WX�0e���Q�j`�����4�.&�:�*��n�e�]�]�*�O`�0�SyM�"�ٴS5�0�NAH&A;�A���W0ΥQ{j�jb���I~m���>�����M�'�K�>����*��~�k~th��U���𶺐�ab��6��T��0�͌X�*��4�����O��ȫb��'[�K����Cي�ž�@���i�C��}RbN�n��VM�B�8�@h�d�ݢx�0)ל"�[(���\-��h���q�G 텪�����'}���^�Mr(���a�}B��e�/?�h����}���B<�S��өS�d2��3a��bʛ`@����5�x{����j�7�Dn�ym��Mֳ������Dn1.���^7��?�Ȓ�`yH ��0y�����0я���j�ֲ�A�dϯ��C:�[�W�"s����@T�������DJ
�+���Y��QW����~�QZ�t���������ċV�?��Vh����A��>��j�����s���;�:g��qK�A�w��[����K$�h�M��������m(�GTY5V���>ٰk{|�tS��v��9�Q��v��4�Y!��a[����A% ����]*x�{\��IR��A�t*�a��k(��A�|�*_K�B(0z!yz�%�^������~��Z*R�5��XL���Ho��?d�`�	�}��L�� �7�,�rh����8J���M�r>r+��(-���ALm���Y��'�=:IhQlv�T��Ȳ;/�'��,^�aDW i"Q�u!5�`�v�Ԣ�;�
�ߙe�ɘ7�� V��{jJ��?�w��vG0�Kxf{W����8�N��+~��@u�-����Bb�����EyTN).���B��˗�f�<�<�힇x�w�˥�H�%�e��s���-���y�G�Ϋ�0��W�}rSǩ�����?B�-=�����-l����y����%���R`����"�2�+W�5��q�.�䘨�Te�D���sɚA�x�Y�o,C@kZ7�!9sV����1��J���U�B��?�Y��Ny3R�:JZ�8�g`J��>��ل�v�r������3
��0f��9�����p��z1�+�c�^�n�]��DkQ}R�vP�75�ܙ'C�'W����3�D��.7�-5�2�Kl,N��IS���*�6��v�h�/�)D?|�.��f �_hxt���}���{qV���{�����s����
�0߻�sG*k����1\4�
�5��:���mDBӆ�0�DcVpEV1MD* TS�sw���Mk2��û �mږ{aO�NҤ-������I�Y�H��56���I�V�Mhl����Š��D�;�������@8��φg�N�\�-�]y ����RNޭ^�����,�ʗ�r�J+�NTᒓ<�
֤�Rg�\�f�H����6gq�A�������7W�p.���#�э��e$���/����k��W���������=�1M��C�<�(_�$��=�c+��>�y�0 b��:8�?ӗ�Uw�ĔK:��C�<�z����yQ�>T}�E�1)�mk��x�����9`����c�cP�kU���Y�	��k��"�tov��
�l#����6F}�6ߤ�K�ۀ�>�H�x>C�=�ߎ=��vk�qU.T�ep�QU�$�Znǉ�O"��f���YYJ��N=��M!��@{�1�#���Y�~���a�F�:�I�pBcD�o��E
�V�:9Z)������ĀW��h��w��l,v`f1n3O�3��lC�n,��5��1��-{d���� _Jx���~��P;J�T�gi��gc�+�
�O�z����kjrZ�g>�כ�aj�����m�z����cj��rdY����O������ki�����8�ԧ�q���]
x�9ԭϮ����v��߭o��{�RO7���K@�ҍ����@��[��8
����i�/�ǣ��������������n���/�'�q��Þ�7A=�n�Nr�{��ܱ#Ѹ�F��t`V�lF��F�1֏4������mj�a�ot�aj�|��H����~Ÿc���zz��|�N��Ξq����ׄ����(A�ǩ�_�Ǖ�����%��b-��3�s
~����v�?D�w�/.቞~��|MC?���ăX.���������K�_�,?�|�]�e��o`�����Ƈ�oż�)��E"�z5�:ʾ]9>=<@~?J^����,��ˮ0z������K=�p�a�V�.uR4�ٞ�����9���HrƸ�T̻���DߏY��ɭ8�vIĕlF��B �k[���o��HϜ�?=�y߇VO��5�� Ƨy����������.��D�mD"�u`q�&��Q�ZY����7
����j��_c�$�Z⸌ �T�i�Г���ch|sGh۲�A�`%�|�9m�϶��I�$>�vw�M�Dӕ:�BX�s��+���*ÆLh�>��NQ:r}g���T����>x�U�I6K�Az�����$�~��k��bF�Xl4t�H��?ږW3E\�N����T;PZ�0L�l�{���4%_�ћ�H<���F,R@�[43:���:j�BnOp���F��7���|�p��5c]�yÏW,+!�-Pj�g����l��7���s�Vj������wk留�m���w���w,x���|��bg
��T�ɞ)�b&�zn��01��_^2g�3*����PwQX� 7�pф�!ʫ��;O��	9xH�P�E���7�9:�X��v�xyl�#��:(Ԩ�d+��.}���
|-������`�j�Q������U�Kt�}����u�d�Y�[`fbK3��D�D���pt�r#����G7h��@�eΖO7���c:0d?w�K�A���a�z@��h�R��q�g`�v�k>�	�wY�󷢾��Ӷ6.��M�Bo��X�����T331���䱟/+�)s�"���`��}��ޢSN�t�g�N��wפ�F��6�s�ǒ�}�f�j���6��l��-�8���N�-�-�!����Չ;x�R�����k�[��i�� b�nh�H�Q�� ����*N�^:����A2�5&ہB-��g�v�5w��t	���,�zD�T��U��l��K��Xb�צ�h��5���o d�s����fV�ݰ�B賢*u��e�����sP .H�`'���.�ܝ����kdK���6�/M\m,��hʂ��5 *���ۼ�X����	�d:�|�c������:��1�"�LU|��Q��L�ǘ��]2!N��%%7�o
Ў��\�j�֝e��|Br�a���9�e�9�]ϴ{I���O����G���h-�C$�nw.~d�x���km-��졘֧��qVu�T�m!�\qp��e��V�a�o�>�OeϤ$(n6��7�F
t�S�y���G7|X�ō,��^\��!g���l���兔������|T%0~��i���Ya�J R9�����(�N�}����}>q��KocG���hBκq��"?�F�Evb��(��C}��������i�0�F�S*b�pW�!`4�Ǖ�me�7{Y�ia;Ny�����ǚ�G)�7K��t��7��pG9��ϣ��Q�ɯ�zUڿQgz�1�a�S�B����'Mʀc�� !u�E���Ɛ��a�%RF�Q�[�Q��x�����5��%�@0u)����A�5�3}��4Oe�P��C��U���D�Ђ��l[p�Wֵ>z!�n��G
�@`lO�����N���3s
�� �l(�i$۽XdP,b�L��-�ˈ�љ�҅|( 3	.��N�}�� �������u ���&;�-E�����,H.쁪8��z�^�Z�=$01}A��ZjC�u��O�Gx�T�k�iC���ay�P��<��S��hΪ"=�bԼR�R+K	FѤ]9�f��H6�q�$ڒ����}�p�uO�5*�qY�r�*6���������]NĈ;�뱩NɷH���T!��R^��������C�`��
���fWE�!������s��,c
�<�T6��I�(�y!��u�v�oZ�=� 0�L��s���gk�w�6�N)m�;���:(�P���R�:*����mQ	V���#�3��d�@l(����dU�ӸJK��CN�+�ϩ���J>�i<����d��u �-�P'g�<���C�:k������"�}���7&ٻ�vU8�b�
%�\5d�_�0|�5Y�X���ڊ�92ư�G�h!��^@,�8��by.e�v�v���d���8��٨�+!в�[t�2�z�t�9q�ZJ��Ft;�E6��8�lх�t����
j�Frv�t{�`��	�z&J��ba�?�tE�K�||�g9�A�CZ���H,r��� ���U|��q:�S뗛%�owI陧���Dã�{�qm�"Gi����]j�s��O��(V f�=���tR�t�2�^-r��d�k��6�+$+���ڣD>�98%�q�Ϟ�Y2�z@�bA62a:���kԉ{ �=2��R`_-��s{N����7�<G=���9�WD��ȍ0������\�9�-~W{F3s�*���٩u�BA�����уq�IA�6Ķ� ג�>�*�U`;�,���1�\v�T��T�VY��-J@;1'�Gf��Ƈd��T����5�V���Pe��y$�vu��E�S�u�ٹ@������XC+4��儃E�&��eQQ�?]�N��)��Jt�.�!i��x��� U�BE�@X�*�����6��[RG�'⛶݆r'��V^������"��knk��g�g��^�P8�v:�,�2���Q�R�^�|�4JA�3�P�M��#]�c��ަCQ#�Y�ai��*,f���[2�	�j�`�Ɓ���gQ��	�k�V�`���mə������b�;�Sq*n�طp�S(͇�=�^ר?�3i��u�s��i�!�H��8H�s����en!ٙ���M�{���J�_��3�)6�,�ń�X �C�k��(=4U4	@q@���4[|.zե~[��E��\A��1ϵ�~���ss�y � p���F��Fn��T�Q��k�J�a�P0�'[6uoj�n�S�;`tP�J��ӂ�.�+X}_˷}�{���� �#�y�2�n�� ��\�j�U���3T�P�c�����M.��({��P�7w�&����km����Ҙޣ���/��I��tz���<YBgf��}��X�\� u>� >U(v�e�ĺn����n����v�ѴF:��cZ�8� 9;��fKY!�]� @����i2q�W>��9���[i����͝��5F�k?t�}>b���I����3�뷛�������1 ������ �,�O/i\���ɸ�@<+>�{��u�Cx��Wp:�� �����`0��o�/3��<����+��W/���7�P-�{&_�׹W��(��O�o���Z&�_�&[��9���'^��2
�/��J?N�꼋�V��ϟ��r�1�������A�+����r�w�s�a���7�W �zb�|�������g��]���=��;��7�\�Y�仺1S` �$@��42`Ѵq߽}����_x����ᦏ�ܬ�ɳ9��}N?l�ǲ�<_x�'����T��2��/�Y��s����l0����%��ݻ�߽���o���9��8 I��ջY�_{���w�O/��ߖ�?��c�}9@u]�_>����g�?�ϴp���v19?. 9?Ύ23���o<���o����O?�?���_��>���;`r������o2���pO�ź ?�_A��?���#�g;�G;��;�ｻ�?��;=�T�8 HᯎM]�~,�	c]���W��ޥ'W� p�\Ҹ� Xs3��R�@���3Zj@�^ ���\����KY=�I��KCƧȑ��@�<qu	&H�V3Z1ثQ��;��gBr��^��j\�J�쪏*�	���R�+1�8�,2������
o�������v3>Tm/Y6gs�|�=#���v"��Gk��� /ݡ'H�;D�T�s����&'ye��T�� [E��2�."(M�x�#]͟��$�6s+J�#�*�&�ӗ�)u��탋
��9'X}]L!��r���������~눗��zU�I����Oa�Q�QU�� ��n0y�}�V���y�E�S��������8!P?/D�Z��lCT?�RE��p3��J��2�򼊙l�~Iok\ZPݫ��Vt�4��m��&�&��
{��M�����j|a��璝b��!�q��`a�� ����6�U��XR�}�%�<��|���F4�o��qtk872�r|��E��P�1+�=H��k:��԰���Cj%�j A��	� .�	[Δ� V�Zy�c��������Ld����8���:W�(+�˪2`�s�I5� Д��Vp����)}(,�s�:�����A3H�w�S;�����o��{?�eՖ9
�+��k1����L�|*9'��8�=dn�����C0���ah$a����ꃒ�V�6DVw�DQ�ˈL����y?kڣ ��H��W�q;_�f���zz{���,����M������>_N��B�z'�G'������x�dƵo�j��<����/�ܽ��2 ^��y���J�;�#�9�W���3`i5,�=���2v�Xp�/�
����u�?��.��D�'�o����ᶖ7��I�J���-�pbXU@r�4�,����upj'�L!jmt!Kw�s)�Ǌ�`ư|I��0 Fgd�3����ӱ
Ļ�CQ��'��I���	[g�IѸ7F�7&�$
��[|4f9�,/h��R��Z.��*>�z
L{B
/���s$n�!�P:�P��C�8s���\[�d�sy.n���hd/9/��� Cҽ5��@bA��	%G��WQ��v����	3V9c��aE�ᦌ��b�d�������v�=|O��ݖ�n���!�G�@홼+V�&��EEf�h4�9�Xf�rt�S!V<����`�!�F��&�[� kwځr����H#40g�������v8��A-��:I;�fzɮ�O�B^�q��W]�w��S�㷰�

e.�]"�:��j�%J\���i��p![qt`%3m�L8=�n:P���ӏ崜��V�6d���s����k9NQ	v�z�@�鑒F�2I�L�ؙ�fj8 ��
�T��E�c��������=���Ԫ�Q�&�,����r�o��/�Pb���=��wQ&F�<A�/VE��H:m�Onk��:�7[\��DEd�>�����XA��ibN�����ߤ�V��d|r��`���@�t#rY�|�[������2�Vc�ȿ�~&E�aÑA�[2~�Yk�NQ�ӿ��{�t7�s�BjŞ�k�Ŝ�}N'^��Խ���C�e^/u�-���4����w#_�,�����ID����GU�޲?tq(LE~&X_�)3�R6o�wM:ڏ��Mr���L���.��ĀM�	i�<�\y�7m��>�xB���e�5���m{�Z=��#�RW|7g]ظrv��3�V�N?2���R\O�+�g
<0F&�˶A�5MZJX8��Eml��Ɍa;,m����U(=���g'y� �����զ�\��v�A��lxQF�y�y���mLb�[��o8�xE�kJ�G�4������_jhp%EuCPY�;�X@r�p�����ȉ��7��Cr��'$�(�rz�oo��}�a���l�u���&�0����#r��O��!ŜT���m�t�ί�O���݆_�>N�7"L,	L	�JM��nc��`=�����߀ɄP�i�ٸFds��"(\!�QMC�>�FW�W'�'k/%����6�^^�P���f[���>�(��������H��cA�Fw�4��������,X���y��ㆺ��A|E�qX;�fĊG@J��Y>��N�f���^7Z�Ӄsk���L;��Ma��'�9iadε<x`�*0��{���5��G�y�/n�8��������Q}SQ6�	�3�3�Bx���ט��4��Cd;�ȍ[�ٶ�y�#${��Wa��hB�e�����&�]U�+R�*�OWq&�W�nGl/�`�gVxL�d��&L����yx����kt�љ�x�:�*�G��X--	.3�[�^��YB(����9�2�~�tǭ~��J�Sfd����x�|����k�|JD�r`,;V4k�S v�u��x�������[{��PR�%%(�r���.α]�M|��O���B��J�+���bE��,�,{c��L�*+��Ů��l�8v��������T�BB��x�J_P�c��tiF:�x�fP����<T��M�Dn.Z���>c��v �v5����"(D�c�.&B#h$�O��\�����ud�Z`dP����P��f.s��x6�7�.h�"��7k�b#�0���l�I'8~q�D�e	�����oI��b��S�N >U��i~�!lg�K��>0��{�4f�ȓItBHUK���z�d�d��X�:G��σ���6�Su<�7��˽l�|���ܯ����,X�(Ȟ�x������;����N�J�o�zG=b�/\����KB�3�?�l��?E�o�Z�C t�3~���/ҥ��;�J�ɊBy�s�A �~�Ԧ������������[����B=��D�-��BK��{xi�w��ciR(O9
�<�)��d��J�=�!~-���dAY��m@"$�S�k��,��H4��; O�v�ÓPm[�Rε��aҵ16f�ۡ���8��f��,#��Fũ�<e��J<E5�TS6?Z��i�:�E��/?N��U���d�aÐ�K��q��%ֆ�[���<p��ɦl*�J�τ�\�}���ˡf�fe�W;B��a-dl����nI
#�dԟ~�X3m��<O<��<�儜�=<ӧ����֒a�p(/qu��Bh�\�	��}�`��zSl��]���y�IK�Q*�M����ʛ�(@m�U&J�/c���l��Z_�śi�L�k���S_�P9����},����Щ��7Jdt�2*_|��M@)\��]��Nv$�I+��.٢E�%�;jz��x�!Y�
	9��u�7}
�.�{aL�� �9��������V��y��ǳ�(�E��D���͘ ��b:�JS��8�9a�̕	���d��+���$��m)�F+i�خ����,J�!{^V9�Z�/̆�r(�o������ƹh�7Z6d�}��������_��~�fq����q��Z��b7�%�C���Qc�9m��pw��AZ��0�Eh^��vZ�)}�W_yP�#�?|/��;�-��ܸ��lnk�.
��l#�J��Qc������A�g���)K}�	�D�Es((=�km�ۚ���H���-�a���T_����8�����X�	(�1�S�@�q�ӌ_L @�>̼����3ű:�oq%Fbe�{�m*�dr�.f�q{�$�ԃ��0*=�$=(3<Q��,x���$ 2���!zX�"o^W��p�̓1�Ku'��P7�CSp�U�}\�}��_�Y���!��'���O[��NI�wOA��p�������+!�;��Ήæ���"��[+ͫ�������F0�q�?�Y�NR�psտop0D��r%	���EE�Ҧgb�o_g{M%)�|<���O!or��Ӷ/T5��`�ãD���ǩ�f��߱��܀}]�v�Co��f���^�4�F~Ψ��Y�����m�� �;^��Ud�e /d4�]�1�5r��-��y�@�� {��� s�~B�'2O�*�}\�c���Hz�|;CE�J��e�U͍/�l�l���_�	����Gڈ�r=.*I�b�.�.���4�(� {�+BW����]2.����z0@Bt>1^G/��:�G�X5�z���8sHG��ݯ+ܥ��)�Uy��16T���P;\ʛ�>U�$0@�T~cA�s8T(�t��k��J~f�"�_-1#ҽ���+�1y�FA�;w��н��TV�u; �(v����DNJ�V�߸�ug���u��(pQ �����rn���׼
d�zUS���`۵1������v"C�6[\%�8Еh����M�aW8*���"v��'�ut�8�1YX��[���Z���V��ZeA� vW��M#�ϸ�Wٲ)i�My�kV*�9�,�F��G�}�1C�{�>6]|���2\�
/x����rݒ�u��g_U���S�M8A���9��@?/h	Ь��p��>�}ź3���m$M+���9g�o�P�� (I�*�|j��@_��~�'���o0 �0>&�P&�[Ħm�Ho�n�n]��ʏ�+�w�L�(j�Y����l.��m1+��BkEկ�����v��.e�<1��ߌ�'ι@��]m�ؑN��e��D�
^�����.�M�b+��<w��0�%2�P8eȝ�� >ԵQ4Ńc�0�'�=�����𕬋x�4��%���������.�n
�����hi�ő�)k���\��i'#���+�*ME���E=����,���oE�os�-nL�MQ�\b�J_+w���N��C�^���~fg��qN��x �W9�����]�Q��_��W�w�������W�<j�Hb�D���#��vt�1+��176X�bh���|��h�d���{��(� q۝��Xh�04���c����n#Hq�A6�W�JBN�����.�cGqs�N$��r�2Oև?&�f$f�p���ۉ�`�D��� ��؄�Ւ)�h��pc�������({���r%����Q]Pb�i�Q�03���r�s��~G���O"��U�^�nx��y�u��]6��C��������b� �GUZ�����5j���_,H�Ԕ����'U�_�*���~��_�Ӣ���;����L�e�Ɗ�y�{�w/,O�d���S\b�S,޼"��~�>��l[�C�Lno���e�E�Lq�һ����f��6�	=��R�o�?���]�zQ�#��З����-���s9�z����O�vV}S/�d�CI7�.���S�o�����19bD��#}	������Rw|���
KR���|m���ӐD��R�MɆ��^ �"�ہ@���<6$�]tk�W�И;<H*��&����-�M������>�(�;�)��;t�2�d������������q�'tX�׌L���Ch��k�B�	u ���x���R�diSͷf�72�u�'4��{&4�����s=>@k3�?��=�1��]�,���;X�'���{/����*3_����"��7���3߹'��7ֿ�7����I�2��<O߄�%�����_�ӷļ��G3ߺ���,��7�O��e��ލ�\�0���Nߩ�0y��M�^35���7�C�O_������f�̚�ʽfl,���^����K���y�"�C�ީ5�3}Um|ť��M�N�ԙ¿�@�ހ��~^��"^C�®~�r�	n%�ī}��A{D�������y��NB�!���5�)��N(�eo>ۏ�뜲/�'�0���o��N]~�3�8��ģ�NB�>���]2�3�4�ݐy��g��b��������a��+�
Ounrqwu����'=��u͊����S6�Ϭ	��_�w3�#&��\��f�"�1&�}�� >S���L�8zL�~z�jj�aUjM�W���H6�	۠*1�b��r��É�0��"��K��ǡ�.�g���ȋ�I�&�ox�s��3�  ��e|�CTp����
�\���z���|84�}0���t��өS&����y_�m��w4�������aÀpb|��cdX��G�I�*>���	/�ȱ�X;U.�Qz����	�|�����[���M�ח$�ỽ�:8%���eu��}+d�@��U��m�o�{��gҩщ��(�y��j����/�n�R@XJ���=���w�|G��vO�K/�@���&���㪃^�~��>m̿6��X,0�Dl�z	�DK�@����m[y}r|���@=��sz˖��z�pur4ɎjGz�h\�t���!�� �<�$v�+7��{}ޞ��\��N��Y�ɷϫ���Aϓ{��n�.g),�ef������������K��kQ,^E08*�-c%<r@�!C����D�-�.�fl�6����;i�p-��'��qȀ�ދ�,�Q�oUP������M�'�����ڛt#���Avn�́D�J-�"��Bӡ���i��ܒ�ǃW��6~
^�
��Ŭ}*��A=�X�U[9���ㅙX�J�ۈ=�d�Rb�j���Γ��>k���e�QݰM���}<Vz������㚤RUaB��W:n�wĊ�v���<���dJ�y�e;k����{��]�@��-��ٖ�:�^�HY��Řc@Lʃ����-1mCo�nֈC����W`�&�Gs:1$b>��1�l� dc�z���S��M3�\�Y�0c�� �h�m�S���Z"?P�y$h�Ύq�Q��������e��!"#«2��%�@�B��X�H"�ji�)��� �v_�"�SR��"*�J��H[���^�g�G��^�aR��V��8ݘW��t�}\�)Gp[:j-Vy=.��f�H�� �s�?!�WE�^����T�f����D)|���2�yyc.�d��H���?Y$i���&N��ݰ�E���2�n���gG�0��J��S���r���
Yf��"'�Ò
~����?"R3A�f�e7��f��d�R��^�P��%=�Z�o\E���q,}rƒ���y�[}����zU�\�&8�!^�v�m�R	b:A�G/(�Ǹ��
��N,3w���B��721���t+��Z<��=\3��qie��Q��5œ��%����E��,QF2�#1���"���}�Q�zd�FHM;�8�ԛ�Q�-����3�D��"� ��~8�¶�X8H�áG�Z�}�����&�������w])�k�E-�yڡA�.L#��}�9�Lk��, ��ܹ&��E4�`Ņ���*j_��}N	�#Ei�WK�7i+��I��땓���� ͐Z�.�� %.r�h`��݊^!����v��A��{zؾ�t�w��a�ω:0S;۳�\��wz���TYa<��\b�2���������|�s�p�Bu=x�,�%
xsc:;XseZ:~��%��sMP?p��XQ��# �2m���m��;tP5�BP���H�k�U#��i��ɑeഷ��5�3J�DCq$���J̟�ϖ��wby飂`���Y�OXjGzq�����81ER$dx����mU+8n�q�^�6��-�/ ��Uk MW,��!9#��~c�Ĉ3�7���.���K�I2�|��TC�I���N�q�u�QI��mi�&�Y#�.�;��w/�5�	�TE�5�qnp�_V�֨�A^����~	�e�>�e[���~4In͇�XA�~y�r�]�~";$��(��וv�S����f�;� ~'����i��Juޜ����@���Tc-}Kj�,��ɒ�iޝe�>.۬�t�FO�	���?}�_�g&��z��z�E�*�͞��i{�G��-�@s���v@'0dAh��]��nݞ΍��`�����u��O�E-ͅ����o��'��n��X����˰������������o��k~��M�����k��W`o��Wj�z/D����I^����)-'���*�����w�7���b���w�&��mŅ�c����k/�n�O~��E�i9� ��-���$^RfCqL�_ޜ�`�{u4��������6�O�cb��ϸ�C�x��>Sy�d����:
x�j�{#�PU�_�˭oV�;�F�r��]�7���oe�����9��=��?}����?m��1��?�6������;����_�ó��;sx�S��O�둙�b�_J-��U[_�?6�������,>Ⱥo=_?�s�A4���:�'�����:��P���_�