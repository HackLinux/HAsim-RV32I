U��j�h0�' d�    Pd�%    Q���   SVW�e���4����E�����}� v�E܉�0����
ǅ0���   ��0���;Ms��4��������  ��4����z uǅ,���    ���4�����4����P+Q����,�����,���;E��  �M��Q�q ���E��E�    �U�RQ�ĉe�E���4����Q�U��E��M��Q�ԉe��U���4����H�M��U��E����4����� ��M�Q��f ��j j ��� �E�������4����z uǅ(���    ���4�����4����P+Q����(�����(����E苍4����y ��   ��4����B��D�����4����Q��@�����D�����L�����@�����H�����V�����W�����H�����P������P�������P�����P���;�L���t�ዅ4�����4����P+Q����<�����4����H��8�����8���R��e ���E�M�A��4����P�M�U�J��4����A��4����E�B�M�d�    _^[��]� ���U���D�MċEăx u	�E�    ��MċUċA+B���E��Măy u	�E�    ��UċEċJ+H���M��U�;U�sC�EċH�M�U�U��E��E��M�Q�U�R�EPj�M�Q�
  ���   ��E�MĉA�%�URQ�e�EċH�M�U�E��M�Q�M��   ��]� �����������U���,�M܋E܃x u	�E�    ��M܋U܋A+B���E؃}� u	�E�    ��M܋Q�U�E�E��M+M����MԋUԉU��EPjQ�e�M�U��M���   �E܋H�M�U�U��E��M��A�U��E�M���E��]� ���������������U����M��E��@    �M��A    �U��B    �} u2��b�E�����}� v�E��E���E�   �M�;Ms
�M��3����2�U��R��m ���M��A�U��E��H�J�U��B�M�H�E��P���]� �������U��j�hИ' d�    Pd�%    Q��D  SVW�e��������Ef�f�M싕�����z uǅ����    ��������������P+Q���������������E�} u�  �E�����}� v�M��������
ǅ����   �������z uǅ����    ��������������P+Q��������������+�����;Es�����������  �������y uǅ����    ��������������J+H��������������U9U���  ǅD��������D��� v��D����������
ǅ����   �M��鋕����+�;U�sǅ����    ��E���M�ȉ������������U苅�����x uǅ����    ��������������A+B��������������M9M�s>�������z uǅ����    ��������������P+Q��������������E�E�M���Q�k ���E��U��U��E�    �E�PQ�̉e؉�@�����@����E�Q�̉eԉ�8����������B��<�����8�����<������������ �������������E�M䉍 �����&�����'�����'���P������Q�U�R�EP�� ���Q�Y  ���U�E�P�M�U�RQ�ĉeЉ�����������Q����������������Q�ԉẻ����������M��������K� �`�U䉕�����E��������������������������������������������������;�����t��U�R�` ��j j �� �E������������x uǅ����    ��������������A+B���������M������M�������z ��   �������H�������������B���������������������������������������������������������������������������;�����t�ው�����������A+B���������������Q������������P�_ ���M�U��J�������A�U�E��P�������J�������M��H�L  �������B�������������MȋU�+U��;U�  �E�M�ARQ�ĉeĉ������������Q�������������������Q�ԉe��������������M��������:� �E�   �������B�������������M��U�+U���E+������������Q������������������������������������R������P�M�Q������R������P�l  ���r�������Q�E�B�������������������E�M�A���������������������������������������������������;�����t��j j �m� �E������������Q�E�B�������J�������H�������������U���t����������M��U�+щ��������������������x�����|�����|����M����x�������x�����x���+�t������@�����A�х�t��x���f�M�f����  �������B��p�����p����M܋������BPQ�̉e���l�����l����E܉Q�̉e���d����U��E�+�h�����d�����h������������ �������������������H��������8�����8����M܉��������0����E���M�+ȉ�4�����0�����4������������,�����,����E��������+���������������������������� �����������������������������������������������+� ������B�����@�ȅ�t>�� ������� ����� ���������������������������������f�f�
뢋������U��������������M�U�J��������������������������������������U����������������������+��������A�����B��t������f�U�f��M�d�    _^[��]� ���������U��j�h�6' d�    Pd�%    Q��SVW�e��E�E��E�    ��M���M�U���U�} v)�E�E�}� t�M�Uf�f��M�M���E�    ���	�U���U�E�;Et��j j �� �E������M�d�    _^[��]�������U��j�h�X' d�    Pd�%    Q��SVW�e��E�E��E�    ��M���M�U���U�E+E���@�����A�х�t/�E�E�M�M�}� t�U�E�f�f�
�U�U���E�    ���	�E���E�M�;Mt��j j �� �E������E�M�d�    _^[��]����������U��Q�M��E�� �n+ ��]�������������U��Q�M��E�� �n+ �M����t�U�R�X ���E���]� �U����M��E��H��M��E���]��������U��Q�M��E��M�H���]� ����������U��Q�M��E��@���]����������������U��Q�M��E�� D'( �M����t�U���R�X ���E�����]� �����������U��j�h�X' d�    Pd�%    ���M��E�    �} t+�E�� �n+ �M����M�U��D'( �E�    �E����E��E�    �}� t+�M���n+ �U����U�E�� D'( �E�   �M����M��U���H�U��
<+( �E���Q���E���A�M��T��U��B�����E�   �E���Q�E���+( �M���B���M���J�U��D
��E��@ �E������E��M�d�    ��]� ��������U��Q�M���]� ���U��Q�M��E��@����@��]����������U����M��E����E��M��������M��AD'( �U����t�E���P�oV ���E�����]� ����U����M��E����E��M����#����M��AD'( �U����t�E���P�V ���E�����]� ����U��j�h�6' d�    Pd�%    ���M��E�    �} t,�E��@�o+ �M���M�U��D'( �E�    �E����E�j �MQ�M���u
 �E�   �U�� 2( �E�H�Q�E��D\1( �M�Q�B���M�Q�J�U�
�E������E�M�d�    ��]� ��U��Q�M�3���]� �U��Q�M�j�M����E��P��R��]� ��U��Q�M��EP�M����U��B��P��]� U��Q�M��M����~r
 ��]� ��������U����M��E����E��M���������M��AD'( �U����t�E���P�T ���E�����]� ����U��Q�M��EP�M��Q�B�M��Q�J�U��L
�U��D���   P�M��Q�B�M��Q�J�U��L
�U��D�P<��]� �����U��Q�M��EP�M��Q�B�M��Q�J�U��L
�U��D���   P�M��Q�B�M��Q�J�U��L
�U��D�P\��]� �����U��Q�M��E�� �5( ��]�������������U��Q�M��E�� �5( �M����t�U�R�S ���E���]� �U��j�h��' d�    Pd�%    ��\�M�h��3 �E�P�[ �����@X ��t�/h�   h r+ h��+ �M�Q�d[ �����_ P��a ���6i j,�:] ���E��E�    �}� t2�U�R�M��?x���E��E�� �, �E��M���o+ �E� �U�U���E�    �E��E��E������E��M�d�    ��]�����U���0�M�h��3 �E�P��Z �����uW ��t�/h�   h r+ h��+ �M�Q�Z ������^ P��` ���kh �U�R�M��>  h�- �E�P�8� ��]�������������U��j�h��' d�    Pd�%    ��d�M�j �M��x� h�q+ �>U ��Ph�q+ �M��=����E�    �E�P�M���w���E��M���, �E��U���o+ �E�j�M��"� �E�� �o+ �E������E��M�d�    ��]��U��j�hC�' d�    Pd�%    ��P�M�h`�3 �E�P�Y �����@V ��t�/h�   h r+ h�q+ �M�Q�dY �����] P��_ ���6g j,�:[ ���E��E�    �}� t?�U�R�M��?v���E��E�� �, �E��M���o+ �E��U���o+ �E� �E�E���E�    �M��M��E������E��M�d�    ��]��������U���0�M�h`�3 �E�P�X �����eU ��t�/h�   h r+ h�q+ �M�Q�X �����\ P��^ ���[f �U�R�M���  h��- �E�P�(� ��]�������������U��j�h��' d�    Pd�%    ��d�M�j �M��h� h�q+ �.S ��Ph�q+ �M��-~���E�    �E�P�M���u���E��M���, �E��U���o+ �E�j�M��� �E�� �o+ �E������E��M�d�    ��]��U��j�hC�' d�    Pd�%    ��P�M�h�3 �E�P�|W �����0T ��t�/h�   h r+ hXq+ �M�Q�TW �����~[ P�] ���&e j,�*Y ���E��E�    �}� t?�U�R�M��/t���E��E�� �, �E��M���o+ �E��U���o+ �E� �E�E���E�    �M��M��E������E��M�d�    ��]��������U���0�M�h�3 �E�P�V �����US ��t�/h�   h r+ hXq+ �M�Q�yV �����Z P��\ ���Kd �U�R�M���  h\�- �E�P�� ��]�������������U��j�hЃ' d�    Pd�%    ��P�M��EP�M��&s���E�    �M���, �E�   �U���o+ �E������E��M�d�    ��]� ������������U��Q�M��M��   �E����t�M�Q�jM ���E���]� ��U��j�h��' d�    Pd�%    ��P�M��EP�M��r���E�    �M���, �E�   �U���o+ �E�   �E�� �o+ �E������E��M�d�    ��]� ������������U��j�h�' d�    Pd�%    ���M��E�    �E�   �E�   �E������E�� t, �E�   �M��A(    �E�j�M������ �E������M��IK �M�d�    ��]���������������U��j�h��' d�    Pd�%    ��P�M��EP�M��vq���E�    �M���, �E�   �U���o+ �E�   �E�� �o+ �E������E��M�d�    ��]� ������������U��Q�M��M��P� �E����t�M�Q�K ���E���]� ��U��Q�M��M����.   �M���`�  �M���$����E��@�5( �M��A�n+ ��]�U��j�h�+' d�    Pd�%    Q�M��E�    �E������M��  �M�d�    ��]�U����M�E��M��U��U��}� t(�M��R� �   ����t�M�Q��J ���U��U���E�    ��]�U��j�h�}' d�    Pd�%    ��L�M��E�    �} �1  �E�� �n+ �M��A�n+ �U��BP�n+ �E��@T�n+ �M����M�U���n+ �E�    �E����E��E�    �M����M��}� t,�U��BTn+ �E����E�M���n+ �E�   �U��� �U��E�� pn+ �M��Q�B�M��D`n+ �E�   �U����U��E����E܋M���5( �E�   �U����U��E���$�E؋M��9( j�UR�M؃��Ԕ
 �E�   �E�   �E����E�j �M���L�`
  �E�   �M����M�j �M���  �E�   �U���H�U��
o+ �E���Q�E���n+ �M���B�M���n+ �U���H�U��
�n+ �E���Q�E���n+ �M���B���M���J�U��D
��E���Q���E���A�M��T��U���H���U���P�E��L��M���B��$�M���J�U��D
��E������E��M�d�    ��]� ���U��j�h�+' d�    Pd�%    Q�M��E��H��Q�E��D�|o+ �M��Q��B�M��D�po+ �U��B��H�U��D
�`o+ �E��H��Q�E��D�Xo+ �M��Q��B�M��D�Po+ �U��B��H���U��B��P�E��L�M��Q��B���M��Q��J�U��D
�E��H��Q���E��H��A�M��T�U��B��H��$�U��B��P�E��L��E�    �E������M�d�    ��]�����U��Q�M��E��H��Q�E��H��A�M��L��E��T��R��]���U��j�h�j' d�    Pd�%    ���M�j$�GQ ���E��E�    �}� t�M��  �E���E�    �E��E��E������E��M�d�    ��]�������U��j�hi+' d�    Pd�%    ���M��E��@�8( �M��Q��B�M��D�8( �U��B��H�U��D
�8( �E��H��Q���E��H��A�M��T�U��B��H���U��B��P�E��L��E�   �E� �M�����t�U����U���E�    �E������M�d�    ��]�������������U��Q�M��E��H�Q�E��H�A�M��L�E��T��P�M����˪
 ��]��������U��j�h@1' d�    Pd�%    �� VW�M܍E�P�M܋Q�B�M܍T�E܋H�A�M܋D��H�E܋@�@�u܋D��u܋v�v�}܍t7�@�D�T
���R�E؋E؉E��E�    �M���	 �E��E�   �E������M���Qj �U�R��H ���E�E��M�Q�Y ���E��M�d�    _^��]�������U��j�h@1' d�    Pd�%    �� VW�M܍E�P�M܋Q�B�M܍T�E܋H�A�M܋D��H�E܋@�@�u܋D��u܋v�v�}܍t7�@�D�T
���R�E؋E؉E��E�    �M����	 ���E��E�   �E������M���Qj �U�R�H ���E�E��M�Q�<X ���E��M�d�    _^��]����U��Q�M��M����N����E����t�M���Q��C ���E�����]� ���������U��Q�M��M����^  �E����t�M���Q�C ���E�����]� ���������U��j�h�j' d�    Pd�%    ���M�E�� �3( �E�    �M���o+ �U���U�jj@�M��4p
 �E��E�� \8( �E��M��d9( �M�袀	 �E��E������E�M�d�    ��]�������U����M��E����E��M��������M�������M��A�5( �U����t�E���P�B ���E�����]� ���������U��Q�M��E�� �n+ �M����t�U���R�fB ���E�����]� �����������U��Q�M��M��������M���`�c����M���$�h���E��@�5( �M��A�n+ ��]�U��Q�M��M��!   �E����t�M�Q��A ���E���]� ��U��j�h�j' d�    Pd�%    ���M��E�   �E� �E܃��E��E��E��E� �M������E������M���3( �M�d�    ��]�������������U��j�h�|' d�    Pd�%    ��@�M��E�    �} �1  �E�� 4o+ �M��A,o+ �U��BP o+ �E��@To+ �M����M�U���n+ �E�    �E����E��E�    �M����M��}� t,�U��BTn+ �E����E�M���n+ �E�   �U��� �U��E�� pn+ �M��Q�B�M��D`n+ �E�   �U����U��E����E܋M���5( �E�   �U����U��E���$�EԋM��9( jj �Mԃ��&����E�   �E�   �U����U�j j �M���L��  �E�   �E����E�j �M���  �E�   �M���B�M��|o+ �U���H�U��
po+ �E���Q�E��`o+ �M���B�M��Xo+ �U���H�U��
Po+ �E���Q���E���A�M��T��U���H���U���P�E��L��M���B���M���J�U��D
��E���Q��$�E���A�M��T��E������E��M�d�    ��]� ���U��j�hOj' d�    Pd�%    ��(�M��E�    �} tn�E��@�o+ �M��A�o+ �Ũ��U�E�� �5( �E�    �M����M��Ũ��U�E�� 9( jj �M���~����E�   �E�   �M����M��E�    �}� t,�U��Bp+ �Ẽ��E��M���5( �E�   �U����U��E�� �6( �M̋Q�B�M��D�6( �E�   j �M̃��  �E��U���8( �E̋H�Q�E��D�8( �M̋Q�B�M��D�8( �ŰB�H���ŰB�P�Ẻ�M̋Q�B���M̋Q�J�Ủ
�E������E̋M�d�    ��]� ��������U��Q�M��EP�MQ�M����U��B�P��]� ������������U��j�h�i' d�    Pd�%    ��4�M��E�    �} ��   �E��@�o+ �M��A�o+ �} u	�E�    ��U�B�H�U�D
�EċMȃ��M�U���5( �E�    �E����E��} u	�E�    ��M�Q�B�M�T�U�Eȃ��E��M��9( j�U��R�M����q����E�   �E�   �E����E�j �MQ�M��   �E�   �} t�U���U���E�    j �E�P�Mȃ��,  �E��M���8( �UȋB�H�U��D
�8( �EȋH�Q�E��D�8( �MȋQ�B�M��    �UȋB�H�U��
    �E������EȋM�d�    ��]� �������U��j�h�6' d�    Pd�%    ���M��E�    �} tN�E��@p+ �} u	�E�    ��M�Q�B�M�T�U�E���E�M���5( �E�    �U����U��E�� �6( �M�Q�B�M��D�6( �E������E�M�d�    ��]� U��j�hoi' d�    Pd�%    ���M��E�    �} ��   �E�� p+ �} u	�E�    ��M��EB�E؋M܃��M�U���5( �E�    �E����E��} u	�E�    ��M��EB�E�M܃��M��U��9( j�E��P�M����6����E�   �E�   �M����M��U܋�H�U��
,9( �E܋�Q�E��$9( �M܋�B�M��D�    �U܋�H�U��D
�    �E�H�U܈J�E������E܋M�d�    ��]� ���������������U��Q�M��E�� �5( �M����t�U���R�9 ���E�����]� �����������U����M��E����E��M�������M��A�5( �U����t�E���P�?9 ���E�����]� ����U��j�h#|' d�    Pd�%    ��0�M��E�    �} ��   �E�� n+ �M��ADn+ �U��BH�m+ �Eă��E�M���n+ �E�    �U����U��Eă��E�M���5( �E�   �U����U��Eă��E��M��9( jj �M����_����E�   �E�   �U����U�j j �Mă�@������E�   �E����E��Mċ�B�M��Hn+ �Uċ�H�U��
8n+ �Eċ�Q�E��0n+ �Mċ�B�M��(n+ �Uċ�H���Uċ�P�EĉL��Mċ�B���Mċ�J�UĉD
��Eċ�Q���Eċ�A�MĉT��E������EċM�d�    ��]� ���������U��j�hi' d�    Pd�%    ���M��E�    �} tc�E�� p+ �M����M�U���5( �E�    �E����E��M����M�U��9( jj �M��������E�   �E�   �E����E��M���B�M��,9( �U���H�U��
$9( �E���Q���E���A�M��T��U���H���U���P�E��L��E������E��M�d�    ��]� U����M��E����E��M���T�����M�������M��A�5( �U��B�n+ �E����t�M���Q�:6 ���E�����]� ���������������U��j�h�h' d�    Pd�%    ��$�M��E�    �} t,�E��@xn+ �MЃ�0�M�U��D'( �E�    �E����E�j �MQ�M������E�   �U���2( �EЋH�Q�E��D2( �MЋQ�B��,�MЋQ�J�UЉ
j�EP�MЃ��  �E��M��t�M���R
 �E������EЋM�d�    ��]� �������������U��j�h�6' d�    Pd�%    ��<�MċE�E��E�    �M��M��U���M��P�E܋M܉M�U�R�? ���E��E��E��E��M��M��U�U؋E�P�M���M��R�E�EԋMQ�U�R�E�P�MċQ��B�MċQ��J�UčL
��UċD���E��E� �M�Qj �U�R�M8 ���E�EЋM�Q�~H ���E������U��UȋEȉẼ}� tj�M̋�M���E���E�    �E�M�d�    ��]� ����U��Q�M��M����E��P�R�:( ��]�U����M���:( �E��M�Qh�:( �UR��3 ���EE�P�M����U��B�P��]� ��������������U����M��E���0�E��M���0�S����M��A0D'( �U����t�E���0P�_3 ���E���0��]� ����U��j�h�h' d�    Pd�%    �� �M��E�    �} t+�E�� $p+ �M؃��M�U��D'( �E�    �E����E�j �M�������E�   �M؋�B�M���,( �U؋�H���U؋�P�E؉L��M�yr�U�B�E��	�M���MԋU؋EԉB�M�Q�U܋E؋M܉H�U��B    �E������E؋M�d�    ��]� �+I��������������+I����e��������+I����ն�������+I������������+I������������+I��XP
 ��������+I��V
 ��������+I������������+I����O
 �����+I����O
 �����+I��8�����������+I�������������+I��������������+I�������������+I�������������+I��H�����������+I�������������+I��H�����������+I�騗 ��������+I�������������+I��(R
 ��������+I�������������+I��8�����������+I��x�����������+I�������������+I�������������+I�������������+I���D���������+I���D����������+I���D���������+I��x�����������+I����e��������+I�������������+I��������������+I��������������+I��x�����������+I��8�����������+I�騴����������+I����u��������+I������������+I�������������+I��xM
 ��������+I��M
 ��������+I�������������+I��� �u��������+I��� �E��������+I��� �u��������+I��� �Օ �����+I��� ���������+I��� �UP
 �����+I�������������+I������������U��Q�M��E�P��( ��]������������U��Q�M��M�舳 �E����t�M�Q��. ���E���]� ��U��j�h`6' d�    Pd�%    Q��SVW�e��M��E�    �E��M�U�R��( ���� ��E������M�d�    _^[��]���U����E�E��M��M��}� t(�M��k� �   ����t�E�P�7. ���M��M���E�    ��]������U���VW�} t7j,�78 ���E��}� t�u�   �}��E��E���E�    �M��M���E�    �E�_^��]������������U��Q�M��M���� �E����t�M�Q�- ���E���]� ��U����E�E��M��M��}� t(�M��&� �   ����t�E�P�W- ���M��M���E�    ��]������U��EP�MQ�   ��]������������U��j�h�j' d�    Pd�%    ���} tGj,�$7 ���E��E�    �}� t�EP�M�蚦 �E���E�    �M�M��E������U��U���E�    �E�M�d�    ��]�U��Q�M��M��h �E����t�M�Q�z, ���E���]� ��U���$�M܋M��o  ��]������������U��j�h �' d�    Pd�%    Q���   SVW�e���4����E�I�$	�}� v�E܉�0����
ǅ0���   ��0���;Ms��4����M�����  ��4����z uǅ,���    � ��4�����4����@+A��   ����,�����,���;U��  �Ek�P��5 ���E��E�    �M�QQ�ԉe�U���4����H�M��U��E��Q�̉e��M���4����B�E��M��U����4���迟  ��E�P�0+ ��j j �0z �E�������4����y uǅ(���    �"��4�����4����J+H����   ����(�����(����U苅4����x ��   ��4����Q��D�����4����H��@�����D�����L�����@�����H�����V�����W�����H�����P������P�������P�����P���;�L���t�ዕ4�����4����J+H����   ����<�����4����B��8�����8���Q�* ���Uk��E��4����A�U�k��E��4����A��4����E�B�M�d�    _^[��]� ��������U���D�MċEăx u	�E�    ��MċUċA+B��   ���E��Uăz u	�E�    ��EċMċ@+A��   ���E��U�;U�sD�EċH�M�U�U��E��E��M�Q�U�R�EPj�M�Q�  ���   k��E�MĉA�%�URQ�e�EċH�M�U�E��M�Q�M��4  ��]� ��������������U���$�M܋M��  ��]������������U��j�h�' d�    Pd�%    Q���   SVW�e���4����E�����}� v�E܉�0����
ǅ0���   ��0���;Ms��4����������  ��4����z uǅ,���    � ��4�����4����@+A��   ����,�����,���;U��  �Ek�P�A2 ���E��E�    �M�QQ�ԉe�U���4����H�M��U��E��Q�̉e��M���4����B�E��M��U����4����  ��E�P�' ��j j �v �E�������4����y uǅ(���    �"��4�����4����J+H����   ����(�����(����U苅4����x ��   ��4����Q��D�����4����H��@�����D�����L�����@�����H�����V�����W�����H�����P������P�������P�����P���;�L���t�ዕ4�����4����J+H����   ����<�����4����B��8�����8���Q�& ���Uk��E��4����A�U�k��E��4����A��4����E�B�M�d�    _^[��]� ��������U���D�MċEăx u	�E�    ��MċUċA+B��   ���E��Uăz u	�E�    ��EċMċ@+A��   ���E��U�;U�sD�EċH�M�U�U��E��E��M�Q�U�R�EPj�M�Q��  ���   k��E�MĉA�%�URQ�e�EċH�M�U�E��M�Q�M��  ��]� ��������������U����M�E�x u	�E�    ��M�Q�U��E���M��U�E���E��]� ���U���@�M��E��H�M��U��U��E��x u	�E�    ��M��Q�U�E��M�U�U��E��EȋM��MċU�+U����B�����@�ȅ�t&�UĉU܋Eċ�MċU܉U�E�P�M�Q�M��6 ���UĉU��]����������U���$�M܋M��_; ��]������������U��j�hP6' d�    Pd�%    Q��0SVW�e��M��E�    �E��H�M�U�U�E�E�M�Q�U�R�EP�MQ�U�R�f  ���Ek��M�ȋU��J��M��f  j j ��r �E������M�d�    _^[��]� �����U���,�M܋E܃x u	�E�    ��M܋U܋A+B��   ���E؃}� u	�E�    � �U܋B�E�M�M��E+E���   ���EԋUԉU��EPjQ�e�M�U��M��  �E܋H�M�U�U��E�k��M�ȉM��U�E���E��]� �U��j�h@6' d�    Pd�%    Q��0SVW�e��M��E�    �E��H�M�U�U�E�E�M�Q�U�R�EP�MQ�U�R��  ���Ek��M�ȋU��J��M���   j j �q �E������M�d�    _^[��]� �����U���,�M܋E܃x u	�E�    ��M܋U܋A+B��   ���E؃}� u	�E�    � �U܋B�E�M�M��E+E���   ���EԋUԉU��EPjQ�e�M�U��M��  �E܋H�M�U�U��E�k��M�ȉM��U�E���E��]� �U���$�M܋E܃x tm�M܋Q�U�E܋H�M�U�U�E�E��M��M��U��U��	�E����E��M�;M�t��U܋E܋J+H����   ���E�U܋B�E��M�Q�P! ���U��B    �E��@    �M��A    ��]����������������U����M��E�E��MQ�U��BP�M�Q�M��  �E�j�M���  �U��E��B�M��Q�U�E�M����]� �������������U��� �M��E+E���@�����A�х�t&�E�E�M��U�E�E��M�Q�U�R�M��i2 ���E�M��E��]� ������U��j�h 6' d�    Pd�%    Q��0SVW�e��M��E�    �E��H�M�U�U�E�E�M�Q�U�R�EP�MQ�U�R�  ���E�E�M��A��M���6 j j ��n �E������M�d�    _^[��]� ����������U��j�h��' d�    Pd�%    Q��X  SVW�e��������u�   �}�󥋅�����x uǅ����    � �������������A+B��   ���������������UЃ} u��  ǅt���I�$	��t��� v��t����������
ǅ����   �������y uǅ����    �"�������������J+H����   ��������������+�����;Us�����������M  �������x uǅ����    � �������������A+B��   ��������������U9U���  ǅ,���I�$	��,��� v��,����������
ǅ����   �M��鋕����+�;U�sǅ����    ��E���M�ȉ������������UЋ������x uǅ����    � �������������A+B��   ��������������U9U�sD�������x uǅ����    � �������������A+B��   ��������������U�UЋE�k�P�' ���EȋMȉM��E�    �U�RQ�ĉe���(�����(����U�Q�ĉe��� ����������Q��$����� �����$����������蒑  �������������ŰẺ�������������������R������P�M�Q�UR�����P�  ���Mk��U�щŰE�PQ�̉e��� ����������B������� ���������Q�ĉe��������������U���������  �`�Ẻ������Mȉ��������������������������������������������������;�����t��E�P� ��j j �k �E������������y uǅ����    �"�������������J+H����   ���������U������U�������x ��   �������Q�������������H���������������������������������������������������������������������������;�����t�ዕ������