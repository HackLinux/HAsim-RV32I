��3���*�ts��߮���\a�*�[ڡ\���Z����D>�NTrY# �|
%D�d$'t�ߩ�_�v���+��'���T��]�u��݃����:����k��<�5��|�b_��d��E=�,���t@.`��]��i$��W��J<fX���,��l����1��2�Ě���\�����%e���ƞ��a���Y�����F��� e�Ϫ�W+�G�j?��p&�vԫ8����.t�9 ������:ǖv���m=Ɠw��Ӫ<��p�X�5��?!�p"�f��h����s��c�,�d�V����z�g���Y��xƋv_��
y�7�S]m���X�
�x����+g���l`�b���7��$V��o�f6t]k24�΋ж���`���E���
��_�V풿���x��R�Ncg��A�ZU���/��ϣ�I��ro������
�`������a�G^"DM�����{m�<���|ff�Uͼ��&�P鲣n�x\���Q�kX�k�a���۾�Qa��Ȫ��L��f����w4��@�O�EmOν��ARÇ�y����]���e��Zt��w�-b,���k�(���S��sb������BY����_��Tv$o�0���w�����UK$f���!��_'�����T�7b����c�3�J����}��O�e�+�P1���Z&�㳅��c�4~�8!-�H�̪�釔������'�ݱ�d��B�"��<��m��
�3o�[PWݞ��f��?�uTߊ��b�9 �#���o�%�rw"x�*lB��O��獡Fd��U��C�)��j�(E`S1���n9���p��L�9��{���؝��K��ֽ������$|���2G�O˭���v��E��	p��hrv��5�E�b�xҮPc2����|��fN8�eDߡq��zv�㳭%�4�e��z�D@T�'���y�鶯_B?A��Y�$�co<{��]٬���D�렐��{�A`lv�Dލ���T윌����`��C�D�̤m�F�fcBz�	����R����:���q���"��F��TT�XBE�T\j�5Õ�1����ͬ[F�!��Wg0�d���#b���E@����a���� ���
eD�c�DU�es���Y�dw�����vcr�iRdܐ� �� ���_�Jo�Q��ۧ�������Qd���e�LT��堐���� ����"zb�e��I��D��]�h!���� �������Jp��k�¸�0�&4��\DTfK�ȅ�����n��Cgd"r�2�m"�B�Ǹ��H����>�B��P��Ccf��fc(��I��Ed��/�U��Bm>��Q�ea���� �b>#o�����L.�$?'C6B�����I*4z1��d������9�슊�dp��a�&%[d��gF��C�Uɳ��u����q��E������A����6!��즿����;`����6�It��x�$r��o�V#C��y��R�㖀�ʑ�a���������rf���t������z��$�����B���7Pr��2P%��m&m�/`\E%j٩&w�tEnDaoE$��u���c�d����I�F�T5xB����a��ϊ���u�7�g��L.��h�T���S����p*eC.���Z�㻞�*��1�K9���+5�LN�4{J��4��ZZ��cx-�S�]�f��7��*8��k;�����g��m��4����w��t�k�%�*)��������Ԃ����b�-���R�J�H��u�
�W�����ɗc���
c�W��b8A9��%v���x�i1�~ EAR#�d9��xө������d8�C�ѻ�"�4���Ċ��<�cL_႐9s
���慷�g�`�e�.��y �a���m���A18�o"�D
�b?�닊�c�����%����*DC�($N��[���G���S`���� ��������#y~��n�0�f��t(bċ�T�����*`�����`R�s�~��r�e����!�������&oe?q9�$�V��'�m��(���Jm��e\��k/58?����YZW�)�^��4>$�:�N�.��z�Cy.���\����p��F��&?4?���W��٭a���{�$K�sӺ*�]+�ky+f��WxN�5㎮�y���#~`�P��@���������`�ɕ�`9A+b�Eb ��[�!��[cC�����.!�Eb\��)��4���;��'.p"A�S��֪&�����2��b�b_9��~ #��Ե$Y��Z�ģd���E��3"��S�jgj	Ea��u�L�5UB����"��Im��#��(��̻�e��j������@u��bߵ3]�@uR�����շ[�e2�b�$LR�乧घ�E��勽ई�$<�o�"T'���Ot��!erNe���X�
���o��Hr��&��ĝ�2,c!�Ð�f}b�Qޝ�M��zd2��]�����]c�G8fr_��һ�c�����".���z��O�5d$�[��J��t�`Le1sZ�64��k���傞ѫ+��-f{�%�X��4�����UÐ�'Mbr_��5��C��S�Ż��Ř�N��/
���j	$��fKc'��AJd:t]��3������,��֢�S����AK�=�_��3`ݔ�ߡKd�]��'`�(�2��d��J`�FÊ����Ԭ��g�����`~��}ᦞY���-a��L�10\�T��0P�����K��$Y�R0�T����� C���a!�tU����z¤�Q'�`w�_�͒Ug{���R����c1�O����F�_��5Ya�v6��:,!\�ْ��d�ޤ���td��Ñ�����8}��\���b}�eh��NDC�2k�U~��U5�Q�2a�	b� ��N��F$N% k�	�����o%����w�hc�	b� �ˎ�#H$N% k��$��E�4m�s�3�#��$^��c��5b�k,w�����d�G���$����ͯ�y�65�]�R���J��K��h�d���&S����q��疄"�E\����q�0�/��ͫ�&+G��TU��Z�Z.����J��/�t����fk���5#����C�VE�J�x4�tf��}f��mf����s�~- �������ħ�����]�柴n��޼���j>x8���t͸%��&�������a6�-���z�e�&��խX�f��^CBi$��L�<55I�5&F��<j�\���J�[�B���Cε4>�eYk��Pz稆̵�\�G^��J�%�떂4�d��`���f]�ǳ����`���Se��._��T��-$#t�K���ɥwab�x#p%2�c�%NC�bc����=�(�>�˺�2p��O�d�:��h���*�LGDUK����\�e��^��Icwe���%�_�uaP�(����ս�;'�&�	��� $��l�[���tL0%�s]a�?�̿���f�f����/�� �4��C���+� �f�Vd"��v��ɖ�s�H�d��'8��|!��L���݊\+�@o���v���n�;ro�(x�n���J4cB���*@�yL�Y���K�����"���a��#@�⊖�Ec ��������EX�c�ʌ��u��S5�h��ɩ?��S��/Y� ��s\�Sde��:"���܋���{6sO����Q*`����?�"�I �I%�O�������&����g�Q��ȄR=�a�g�
��x#G4�����ڠ�eC���a� ����dS�KS�ʕaqEd�B? �+�����ʎP�Ͽ�ĵ�mbB4�5�� Ǫ=��d����=�b��dx%��~�@WY��{����e���?7�������=dgaC''4�����xҮRcR�M��|��:oC�H��(A�^Z�"Ї{������[�&�ɽ�by�q���$��.���W�l�Y�˹M����qd�i��ɠ��z��R�8�.��s~$ �N����<�G���,���yŠ5'4���.��9!�۷b5�nPc�F�'�����r%�ۍ��D��*�|#9!ň��7@�C&�����s�����d���b����e,9ҥi�cwd�e:��"�?�"ï������4�E}�pȝ�����e���D���d�����p� ��`�:��Ն|��sƥa� �w��toCtd�3�
�����Pcr��鍃�_ ����|Ԩ�,���-�����<jUb��_�&��Ֆd��4����&@u�č��Y�f0x|��A���`��B:�����b�ry�\�������� �ͨH����[ �̯��w���\�#���"��d�����O��҅���]����gѣ��冇e�s@D֣3��2��?��F��6�c��TςՅ��5��զ�g6�����cWp�A�e�Ǆ���U߯Y�N�Q����囷+���<�i����f��e��?9e�w���	��M�'��bp`V�3l��s�;�R�������5�a���B��e佘'e��_<�/+5F��O���OGb]����U\c`���xMr�J��g��^�}��,p�5$ �������1��W��ѿpP���Ł��uϪ��N�o�l�֙�N��������t8���b
�>�UJ<��Q�S@|�d�`C�w�ρ[����"��W+a���lb�����R���t$�s*� +\�6���/7�CF#>�4�`���\7��#5����2�øG�5f&�k����Qf�R���y��H��=#@���!�V������S���#C�ׯ�'%`�b�bs��B�|���|�G��n�j��G���[��Md�f��ⳮL�A6��������策�:�A�鹌�|��9��%��K�Bȳ�������q����p ��Y��?�T	ϝ9%�Rh��" �+����]�,���2��cYب^&�5;gݥT�(�������H}d�I}coeʢ[e7��%n���﮿^ 6�����c��1���|g�ࠊ��ڙ�k��G�����%�[���K��|�����LЂ=3��~i�С�����1������A00�ߩ��v��o��#���:��@ł����-x�Nv��\����έ2���$F�����i�&B���6�`l�_�����w1�y��ʡ��p��0��LR�� ��1�憞�o��a*��:�����ED����V>ty� @#��G�8!Z�ǿ�����2��:P6pZ
q։ 2��	0���sc�9�}{�\�i�}��h��uY�����T"���"����;�$����q�%�ĂR�K/��(����eĚ�m�:
�~�U�NR�)�D����Z���$�K��`�+�������=rF�MScb꓀w�aS��U*RB8�3�iܬ�d����/�?�ܯ���~!�"פm�N��|�T?�/��E	�5�,e����s��\�UO=OdÓ�Uj����r� ��tvA�u,�� M��r����DO���"U�!��,���R�:�K��#�b�������E��sg�뤦%%�ͤ�������o4��'�ZDa{P�͋[3����,�3��#D�5v廢"YC[D+j��4�U�J�!K�11����+�4g�D?�v廢���3������8��=L��E����L���+�4��6P���Yh#OC[D+j�`7�U�H�)k�Ɏ�n��o%���d)��Ǚ¿�3������H��=L��E���|���+�4g��e.���ʺ1��jl_[��,�lGs�V��4!��7������)�`7_y$!��]^%�Q�c��R��(� 쓕e���֍{�*�7�%��gT�������Ó�r(M2Npps�(��%��E�L���mݦ�*4��ע����J���*5��8~���$��b�Ӄ��4c�ez�,�z�=����2�&��n#o�w�����׼������2