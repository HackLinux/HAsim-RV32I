��������������������M�M������������LLGG>GGG>>5>=/>B??>DBC@?@D?B?@CKB\D@\BDD\�\K��\KDDDB@?==D=>===/=>>D@BLLGKGGjLLLjH�M�����M����������������M����H����k�����������������GG>GGGj�������������������������������������GGGGIG>E>>E/E>@>>G@G>>>GGF@G>LGGGGLGGG���������k�����j��LLGLGBGG�G@GDG@B=@>/>5/>>=/5>/5>GGBG�L������M�������k�M���������LLG�GG@B@DD=>//=,5==-.557-,(.(,*(&,*&'%&&&+(&%&%2.77.777.78...+.+.7.8..6.+6,.+.'.6,+..6.,6.77.8..7....7.�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.>?��������������������//>>>GHGHLLM�GMLGL�}�yddcdddcVVVUQQRQ
-////E>>GGGGGGHLHG�M��M�H�������������M��M��M��H�GGM�LH��LM�M��HL��G����M�kM����������������M�k�M�HGGMLGGLLGGLGG>>>G@E@GGGEGEGLLHLM�����������H����M��k���������L�GGGGG/B>@>>5-/?=B5D?=DB?BC=@BD=C@CDDD=@\\DD�\B�o@DA?=B?5===>==--?B>BDG>KLGLGGLj�GH�M���H�����������������H��M�jM�kkH������������������GGG>GG���������������M������Mk���M������MjGGGGEGG>G>///>>>E>@E@G@G>>>GG>GGLHGLGGH���������������L��LjLG@BGLD@GG@DG@@>5=>5/>5>>//E/@GBGG�G�����M���k�����Mk�������G���LGDGG@>B>>?5-/,5=-.-7(57-.(*(+(%&'&+&%%&%&%%&
7.77..77.7.7....7,.777...++6+,,.+.+6+.,..+..77..7.7.7...�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I8@>��������������������/--EGGGGGLHG��HG�Gl}}ddcVcdVUVVUQURRR--E-///>GG@GGGGGGHL�H�M�M������������M���HM�k����Gk�LHLHG���G�GM�HLHM�����M���������������MM���H��LG�GHGGGFGGL>>>GE@E>>GEGGG>GLLHLHLM���k�����M��M�������M��H���GjGGBG>>>B>>>=/5@===5==BD===BA=?=@B?\D?@DD\DDC@CD�=B?B?===5?5=>=-=>?>>>@BGLGBGGGLGG��j�������������������M�����k���k���������������������GFGGjL��L������M����M�������M����M�M���GGLGGGEG>>>G>E>>>>>/E/G@F@>>GFGEGGGLLLG����������M�����HLLjL�LGGGGGDGB@>GD>>5>/////>/=>>/>GDGG>Gj����M��M���������M������G��jGDGB@B>>=5>==-.55-.-2(57,(*(,&+&&&)&%&&'%
7777778..7.7..7=.8.77.7......6..+.....6.+.77.78..=...8..�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.@@��������������������-(EBGGGGGHL�H��LH>}}lcUUUUUVVVRVQRRRR
---/E/E>GGELGGMGGGM�H��M��k��������k��M�H����H�M���LHLG�GH��G�ML�GHL�M�����M��������������MH�M�Mj��GHGLGGGGGGGEGG>>EE>>>>GG>GGGG�G�G��M���M��k���k���M��M�k�jM��GLLGG>F>>B>/@>5>5=>==5=@?5B?=@==BAB?@DDBDCDDCDBCDD?BC?B57/==5====>/=>B>>GBG>GLG�GGGH���M�M���������������kM�k��L�����H��������������������GGGGG�G��k��������k�M��M�������k��M��GH�GGGE>>GE>>>>>>>>>>>>GG/>GG@>>GGGGLMj��H����M��������LjG��GLjLLGGDG@@B>GB>>@5>5--5>/>>>>@FGGGGGL��������M�M����������������GGLGGB/>5>>5=/=/.5.-,-,2-*,,,(*&%&%&%&'&%&%?7?7=7.8.=88.?.87.?.77.7.7..7.7...7.7.7.78.778.7.8=8=.8.�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.@/��������������������(-->>HGGGHL��M��GElulUVUUUURUVRRRRRRR
---E/>>>GFGGHGGGHLM����������������������Mk���k�M��H���M�GMjLH�GML�H�M��������������������k�k�M�M��HGGGLLGG>GG>>>E>>>>>GGFGG>GGG�G���M����k��M�M��������������jLHGGG>G>>>>B>>==//=?5>==A===?5?=A==@D?DDDD?DDDDDDCB?@?=>=?55=>==>==/>@>@B@BG@GG@GGLjG�������������������M������Mj�M��k����������������������GGGj������M���M������������M��������LLGGGGEG>>GEG>>>E>@>G>>>>GG>FGGG>GG�G��M������������������Lj�LL�jGGDLGZG@>G=>>>/>5//5>>>G>>@>GLj�H��M���M�k����������M�M����LjLG@G@>>>=>5=>5=-.5-.-,-2,,((*('&%&%&)(%&%%%A=87=88=88==8?78.8..7.8...777..78.77.7..877?787=8=8?.?.7�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I,?>��������������������-(->FLGLHGM������-V`VUVSQUQUQRQRQRR`P&
/-/>>>GEGIGGGGHLMG�M������M�������������M�M�M��M���G������GML�LGHLMj���M����M�����������M���M���ML�jLGGHGGLG>G>GE/>>>F>>G>GGGG>�j��M�����ML���k����M�����M����LjLGG>GF@>>>@>=>5>/=>==B?====?-==@=B?DD?DCB@D\DK\BDC@B?=====5=>====>5=@B>G@BGBGG>GGLjL�M������������������M�M��H�j����kk����������������������GGGj�������M�����M���������������k�HLHG@GG>>G>>>@>>>E@>>G>>G>>G>>GGGGL�H����������������M��������LjLLLGjKGGDB>G>>=/>/>5>>B>>>G>GLLj��������������������������M�jLGLG>G>@>5@=/==/=-5.5.5,-.,,*&,+&'*('&)%&%%%%8=8=8=7?8=88.7.=77.8.=..8.7.7.8=...777.7=.8.8=.8=8?.8?88�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.@@��������������������-&/>>GjHLLM��H���-V`RUQQQQQQSOQORRP;R
--//>>GGGGGGM>GHL�����M���������������M����M��M��kM���H�����G�MGLLM����M����������������k�M��k��LG�LHIGGGLLGGG>>G/E>>>>GG>>GGGGGG�H��H����jH��M���k��M�M������L�GGGB>>G>/@B>-=>=5====@==@======?==DB??BCDBCDCDKDB\@A>=7=====>7-==>=?5@>G@GGDGGGFLGLL��HL����������������������M�G���Hk�����������������������GHGj���������H���M�����M�M��M�����LGLGEG@G>>G>E>>>>>>G>G>GG@GGG>GGGLLM�G���M��������������������GL�LLGKGGLDGDB>@>5=>/>/@>>>GG@GGj�������������������������������GGG>@B>>=B//5==/.5.-=.-.2(.*&+(+&'*(%'&%%%%%=7=8==87??77?887.7877777.7.78.7778....8=78.==8=8=8..?..7�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.I/�������������������������HL�HL����M��A[J[\nonronorOORPR`P->E>>G@GGLGGGGHLM����M������������������������k�M���jML������GGHGMLM���H���������������M�M�M��M�GH�GLGGGGGFGG@G/E>>>>B>>GE@GGGGGGG�L���MjLMG�M����L����������GL�L>G>>>@B>>>/>=/=>==/====B?.==-=??=@C=@CBDCB@CBC@?DC===-?==5==/====/>=>>B>@GGBGB>jG�LjML��M������������M��M��jM�LHM�k�H������������������������GGjj��H��HL�H������M������M�M�����GG@>GGIE@G/>GE@>>>>G>G>GG>>GFLG�GH�HL�������������k��k������Lj�L�GLGGDGG@DG>/>/>>@>/B>>B@GDGLLj��M�����M���������������M�����GGB>GB@>>?/5=/=5=-7-..5.-,+(&,*,)&,%&)&'%%8?8=887?=78.8?.87?.777777.7777.7777.8..=8.7888.8=8=8/88.�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I,/@�������������������������Gj�MLH��M�HLAC<[[no[onnor-/>>>>>G>GGGFGGGML�H�M���������������M����M��M��M��k��LHG�HLMGGGLGLH�HLM���M�����������H�M��M�LG�HLLGGGGG>GG>GGE/>>-E/BE>>>>G>GGGGGGHLH�LGH�LHL�MGk��M����LHL�LLGG>FG>>>@>->5>=5/5==-5=====-7=/==C=5=?BC=@ADA@A@?B?====.5=?5-=5==/=5=/>=>B>@@>>G>GG�jGG���������M������LMj�H��Gj�LMk�Hk�������������������������GGGj�LM�GjML����HL�M���jM�L��MLjGGEGEGEG>>>E@>>>>>>>>>G>G>>>G>GG�LGH���������������M�������Lk�L�j�GLL@GGBG@B/5>/>5B>/>>>G>GGGGGL�����Mk�M��������������M���L�LG>G>@>G>55?5==//75,-7-,.-**,&+(+(%&')&%%%%A?7?7..788=8.=77=77=77.77.7.=77.7.7.7.788888.=8=8=8?8.?.�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I,I?�������������������������jH��GH��k�LL8AYJCn[[J[nno	
(-/E@>GEGGGGGGHGLGM�LH�����������������������Mk�M������H�L��G�G�HGHGLMGG�M�����������M�M�Mk��M�HGGGGHGGGGGG>GG>>>>>E//>>//E>>G>FGLGGLHLLHGLjGMG��LGL�H�L�H�HLL�LGLG>G>F>>>=--5/=/5==-==/=5=.==-=7==5.5?=@=B?D=@BC@=?5==7/57=.-,5/=5=/=>/>B>>@>GB@G>LLGGGjLM����M����������MG�MGGGHG��k�H��������������������������GHLjHLLMG�H��M�jH��M������H�LLLGGGG>>@GE//>>>>E>@>>@GF@G>GGGGGGHLGLk���M������������M�����jG��L�GjLGLDGG@G>G/B>/>>=//>>B@BGGLLj�M�������M���M��������������LG�@G>B>@>-5//=/=./5.5.=-2,.(,,*(+(%%&%&'%%%8A=8=8=8.?78=8=7878.8.8.77.7.7.8..8.7777=.7=888?7?=7?.?.�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I,/@.//���������������������ц�Mj��M����H8:[YJ[C[JCC[n&--/E>>E>G>G>LGGLGHLM��H��M��������������������M��M�k�H��LHG�GG�HGLGGGMGLH���M�����M��������G�k�LLGHGGGGF�������������-E-E->E>>>G>@GG>GLGGLHL�GGHLHGLH�G�MjL�GGGHIFGGGB>>>>E=/>5/=//5=5-7=-5=7/=2/7==5====??==A===C5==?==5=2=-5.=-5.=5/=-55@5>>B>G>GBGGGGLj������LM����������L��GG�GLMk�Hk���������������������������GjGGLj��G�GM�G��H���H��GHLMGGGGGG>GEG>>>>E>>>>>>>E>@>GEGG@GGGHLLHLM��������������������������j�LLLGGGKBG>@@>>>5>>5>>>B>G>GLGGL�j�������������������������HLLGGD>>B>>/>5=/=-5=,5.5..-2-2,(+(+&)&'*%%&%%=8?7?78=.8=.877.777777777.87.877.7.77.=77788.?78.8888.?.�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.I/=./���������������������цk�M���M���j7:<A[YC<n[C[n/>E>GE>>/>>/>GE>>GEGGMG��G��M����M������������������M������M�LH�GLGMGGLLGMGGHGLM�M����M��M���k�M����HLLHLLHGGGG>�������������----E-@>>>G>EG>FGGGGG�G�HGLG�G��LHL�GHLGGGLGGGD>G@>5>>/>>55>55./-.-=.5.=5==7-7===A==AB==B=7/A========-257-=/.5=-=/-//>>5>@>GK>GBGLL�Lj���j��L���������jLHLL�LGGk�kk�����������������������������GGGH�LH�LHL��M�LM���GMLGGLGGGLGGG>>>>>FG>>>>>E>>>/G>>GGGGLGGLHL��M�����������������M����������jG�GG>GD>GB@>G=>>>>B@>G>DG@GGGKj��M�������������������M����G�GGG@>B>>=@=>=5=./5,-.5..-2-.,*,(,+&,&%&%%%8=878=8=8.78.?..877=8777.7.77?.=777.77778.78.?8=78/87787�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.@@./@���������������������цM������M��M::A:ACCYCCCCn>>>G>>GE/>>EIF@>EIGGFLGMLGMjM�����������������������������k���M�HGGHGMGHGLHGGMLML��H���M��MGM�M���M�GLHLHGLGGGFG�������������(-(E-E5>E>FFGEG>>GGGGLGL�GGG��H�LG�LG�GG>>GGG>GG>GE=>5>5B/-55-55-,*5-55=5=/.55==========>755=====5==2557=5=5.-55/=-5->5>>@>>GGFGGLL�jLLjLM�jMG�����LM�LjLj�LLLG�k�k������������������������������GjGLLGMjGLH�LM�GLMGHLGGGGGGGGG>G>>GE>@>>>/>>>>>>E>>G>GGGLGGL������M��������������������������LjLGG>GGDG@>@@>>=B@>B@@>GBGGGGGG����������������������k���LLLGGD@>>B@>=@=/==-=.5,-25./,,5,+(,,*,*'%&%%&%??77.8.7.78=887?8.?8.8.8=.87.778.7.7777=.?87.8.8.?8=....�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I./@/=?������>FGGGGGFL��HL�H�����M�������M��GGGHLGLGG>EG>G>>G@>/>>G>>>EIEGGGGGMGLM�����M�M�������������������M��GHL�MjGGGGLGGLGGGGGGHLGM�GGH����LGM��k�HLHGLLHLGGG>>>>�������������-&E(E-EEEEEEFHEE>@GGGG>GGGGGGLLLLGFGLGLGGEG@G>@FFFFFFFFFFE5E-5E55E---5555555->5>5>>5F5=5B5=5-5>F55E55-5E55-F5--E5F/EE-EFFFFFFGFHGLGjLGGG��jLjG�����LLHGLLLjGLLGjHHH�������������������������������GGLGGGGGHLMG��GGF�LGGG>GGGGG>@>>>>>G/>>E//>>>>>/E@GGGFGGGGHL�jM���M�����M���������k�������GjLLLGL>GBG@BB>>>>>>@>@G>5>GDGGG@GL��MM���k�������k����M�jH�LGLGB>>>@=B=>?5-.5==5.-.5=,7,,,*,(,,*(+&%%%%%77777.7?.?7?..8.777=7.7.777777878.878=.88.?.88=..=8.8...�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.@/?/=������>>GGGGGGHL��M�jM��M��M��kMk���HLGMGLGHGEG>G>G>E@E>E>>>E>>EIGGGHG>GGM���M�M�k������M��������M����M���GH�LGGGEMGGGHG>GGGHGGGHGGGGMLHGHGM�MG�jGGGHGGG>GG>E>>�������������E-EEEFFFGFFHHFHEE@>GFLGE@GGGGGFGG>GFGG>>>>GFG/GGHFHEHHFFFHFFFFF>F5FF5BBFBBEB5GBBFBZB>FBGBFBG>BBBBGBEF5GBFB>F>FFFGE>FGFGFHGHHFHHFGGDGLGGGLLjGLG�L�L�LGGGG�GLGGGBHHkH��������������������������������GHDGGFGLGLGGHIGGGGGEGGG>GGGE>>>/>>>E/>/E/>>E5/>>E@>LG>GGG�LMj��M�����������������M�����MLLGHLLBGGG>GBG>>=>5G=B>>@>/>GDGFGGGG�LM���M����k��M����M�HL�GLGGG>>>>@>B//=/.5=/7-.5,-7-7-,,,*.(,&'*%%%%&8=777.78.8=8=8.88.78..7=.8.=77/7.8=.78.7.?....8=88?.....�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.@?//I������G>GGGGGGHLM��M�M������M����M��GHLjHLLLGGF>GGG>>>>E@E>>E/E>>EG@GGGGGH��M��kM����M����������k�����kH�GM�jHGGGGGFGGGGFG>GGGGG>GGGHGLGGGGGGjGMGGGGGGGGG/F>>>>�������������--EEEEFFFEGFHHEE/E/B>G>GE>GGFLGEG>G>G>GE>>>/>>>HHGFHFFHFFFFFFFFFFF5FEFF>F>F>FBFBGBFB5GFB>BF>BF>BFBFF>FBF>FF>E5F>FFFFFFFFGFHGHHkHBLG>G>LjGjGGGGGG�G�GjGGGGGLG>G>kkHj���������������������������������jFGBG>LGHG>GFGGGGGE>F>EG>G>>E/>>/>>-E-/>/E/E/E>/G>GGGFGGML��H�jM�����M���������M��k���kG��GLGG>G@>G>G?>>=/@>G>=>>=G>B@B>G>>�H�LMH�M����k�k��M��LGHGGG>G@B>>5@=B=-=-5=.=-.*-.,5.5,.,*(.*.*'&%%(%'7777.=..77878=.7=.8=77.8.778..8.7?78.=8=8.?.=8=8/8..8.8.�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.@/?/@��6��GGGGL�M����M���M��M�����M���M���M���HLGLFGG>G>GE>>>GG/>GG>G>GGGGGGLML�M���M���M�����������M����M�Mj��M�GLHGGG���������������������������������������������������������������������GFF>>G>>>G>>>G>G>G>G>EGGG>>GG>G>>E>GHF���������������������������������������������������������������������������HHFGDGBGGG�LGj��L�LGLjLLGGLGGjBG>>�kHj����������������������������������GGFGGGBGGG>GGGGG>GGGG>>>GE>>E>>/>>-//>>>>/>>G>F@G>GGGG�G�M������M������������������M��j��L�G�LLGGDBG@B>>G>>@>B>>@G>GBGGDG>�������������������������>>B>>@>>>=B=/=5.>==7====5.57/2-,.2(,,*'&%*%&&%%8=7787.78./8?.8.77877.8.7777.77.7?7.8.87?88..?.?.8=8=.77�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I,/?/=I��.6��GGGG������M����M�������M�������������j��GGGEGG>E>>GG>EGG@GGGGGGHMGMG�M��M��������������������M����jM���GHLLGG���������������������������������������������������������������������FGE>>B>>G>FG>F@GEB>GEG@GF>G>>@G>>>>FFH���������������������������������������������������������������������������HjHBBGD>GLLLGLLj��j�LLjLLBLGGGDG>B�HHG�����������������������������������GGFG>GGGGEGGGG>GGG>LFG>>>@>>>/>>/E-/>>>>>>>@G>GGGGLGGHL����H������������������������M����LjL�G�GGGDGBB>B@>B@>>>GDG>@G@>B>�������������������������=55>?>>==>===-=?=======?====7=.-2,,,*,&)(+%&%%%%%=7?8..8=.778.7=.87..7..777.7=.8.8.78.=.77=777?78.?8.?..7�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I,?>=/?��?C��GGGG������������������������k�����k��L�GGGGGG>GIEG>>@EG>GGGGGMIGGGGM���������M�������������M���M����M�GGLGGGG���������������������������������������������������������������������FFF/FB>E@>>B>>>@G>G>>B>>>>>>FB>>>>/GHE���������������������������������������������������������������������������HHFGBGGDGGGKGjLjL��L��GLGGLG�BGG@GGHjH������������������������������������G>BGGF@G>>GGGEG>G>G@>G@>F>/>/>>/>/E/>//>>E>I>GGG@LGG�LM���M�����������������������������GLjjLLLDGKBG>>D>GB>D@>G@D>@>B==-�������������������������,(5,///@5@=/B7-=?=-====B===?-=7-2-.,*,,%,&)%&%%%78.7.7.?77.?.877.=77..?7778.7777.77.878=78..8.8/87.?.7..�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I.I/==@��@C��GGGG��H��������M������������M�M�����k�GHGGGGLGGGEIEGE>>GEGG>GGGGGGHMLM�M���M�M�����������M�����k��M�LHGGGGEG>���������������������������������������������������������������������EEE--5>/>E/E=>>EG>@>>>>>/E>>>>>5/E-EGF���������������������������������������������������������������������������HjFjB@GGDGGDGGKjLjLLjLGGGBGGLGDLB>kHHj�������������������������������������F@BG>GG>F@>>>>G>>@F>@F>///E>>>/F>-/E//>>>>FG>GG>GGGGM�M��������������������M���������jLGLLGGLGDGG=B@>B@G@BD@>B>B>/==-.,�������������������������)(*,-,/>?=5?/==/=.=====?5?=2-2,7-7,,,*+(%&%%%%%7.7.7.7?8..=8=..8=..8.?8..7..7.7...877.8..7?8..7.=......����������������������������������������������������������������������������������������������������������������������