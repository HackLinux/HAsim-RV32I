�����E�ԓ���6H@Kj[KGu��￁�FcE����)z�
���9�xC�Jm����8|���Yl���%T��x��:W�b�"���=P�.��~��[��:�E2�:��n��Wus���&�f2�KAd��F���'���C�z6#�劅��W�ɢ��$������
�Q��c�����0��!c��#UE�?�j7���g7 ��u�252�CG@�{y�j��=~'P���N&[3S9�
�����E.�a��ý(m�!ǟ��T<�4���\|��U4��`'\@��b>K��) 倇[M�6I�^�{$�V�]UQcd�9�x�P�?�y���uTVj%�ӴC����!�N.��Gwn�H3�ڠ!WŠ!��~�Bqn��")�^�T�}��{�'�LQVj�Z����^�q�ώ���al5Ҩ��+V��r������;�'l�G5���+����b�z�h1OF�C�;����W1=�-��gה��z���0/Zzτ>���	��793�aG�m���E9��&��mJ�=�]��Y`��D���P)8�QWb4/AETfCZ��q��S�Ik�����(��
�����"����w/�%&l)�҆��1bH�����Bv/��TqUH�4�D�:wk�;�~a#.�ń������q��Vڈe{鉘o���'br�a	eZ0/2����Y)q���������.9��G�U�嘉]�R�:�,f��$-����0����c�g��g��~���e�!�|>*�\i�4��m?�G4pj%��_W���-����T�=��F�2�Q��v�!Qk�����qբ���#Q�9�gmF�6C4(���M92O�Q�^�1X�Q3�%�C�)��I�~��Y���C=�+X�� ��"�����#���~��9���8�e{%?���s_!Z�%�V"�����޷��-eE���)��F>�
(!/'e_)��Z��JDB 2�b_�P:��1B��CCCP0c7�Q���qz�5�]B��2����}+�F����)�?���uX����3W��4=�Pz*�v��0R	ۡ�3�0�E�>��>F����޹ ��d�]֛Eu�V�;	��������F�5=�e�گ���}�`�nM����\�*1촋좙7zy#o{SO{;�$|���d��c
��;Œ��x�eQ~��L�z�B� ���A̛�˼Gz�&7�X����'�O�L�t���^'/3�Ѹ/�&�^��<���]Z���{K1�g~2�CgYt����mυe
�)@RU�VJ"+��z
�[H)������*up�7�E�ٰ̎�j~2�n��_�`	ꅕ}-��{�f ���(��u�ň.L5~��?ʞ���{����&S��&�NpJ����4(y���R��:����dyM���b�Ds����K�8�Zt*HkAY��,����{�fe2��u<k�����?�ϒ)�EY-4+y��cU1�4��ʴ����J�������\7����}�Z�k��		t��g�^�����eN��b�V���l�F�I�*��̼��$�i'����3���O4��<ϣCe�₞����/�b�W��x�5����S���]��g��	��¤"Wso�{�/T�`(�g`"��6����0<6� ����/��ó�n������?���d��W���UQd���A��<e��{y������I��{h%�*?��B$�'��5�Ɣ�磱�V.���µ��*��g@4��< �r����&���y}?�/�S��H8ň��Y?t~��"d�Þ��T��EĲ���(i���u�d1�"�'���=MQ������~���m�?�z�~o;[����T���"���D�&����"�"��.�u�\r��|*�k�0F��0��{������#g�ԟ�%~��(�"����P���9T��(�UtX f�:�m��W����B[��:.�<.�n"���] �q>
�S�����0�E��&��R�aQV�i�b�Z� ��?��
���\�XK�D�dZ���Y�hA������}?��>(�5��(��U�Y+�2M�Jb#�\�:�eV��9��"�/��)V���)\��#� �S9�v~��$r��$X�(�F���bS���&S��}�>�M��V��o�T��� ��?����Z�Z��͇
�Pl�协D
l�D*U�1ά�]��"��q-	��m�{��bvd�!M����d%�O�0RKX�A?�7vu��9//ӈ��a��o�\ ����w�j�b�%b���V���-d���^.:�O�����7�4��0�d�Q����Ma������
�GA�b����*<�ɓ����������C�i��%�Nx^�Gyh��sQ������ � �n�w�����'KD\�^����&LNc���n?�Cr�0[��o���-d��B7ԉ�����p���1m���D�7����ECZ����7�O5Psc�v*�����'�4�i>G=�^`2N<���C�	���cSn���+cQ��]D&�pk���Lbk`��JT}a��9۶�&��ͺ����Ŝ�F�5�����^@ܠ����B#�Ы:E��w�S�'��/���ܔ��fs���n�(��u��ä��U &.��k
Ǎ`�����Eq����Âw�)��bu��ab�ףfԷ��Ŏc��f��%����v�Ũ'�׌6	K�J�X�Bմ��#g��e�k�d!�+?�m��U��d�,8�um�H�� ����/����s�&sLꭤ�����`��'f�J¼���9�!:�k��-��E��r���wd?h��D�I$�_I��Mz�G2�7�~\���BVB!h��{��fځ��Le���"ܧ��j߲8�C�
��;}pQ1�q�4bD$�҉F#�lY�d���f�+B�!qr��R����U/�%e���J��H�b�f�ë�S���(x�a�<7��g���}7�c���/TPŁ���'����ѧ��i}�����L��dr�Q�ؔF��z����������������]�tc��f���,&"Ŧɥ�E�S�W��&��F��%̀�e�Օ�V#���ߵ��j~�R=3�-g����k�n~ᶘA�kP!��w{Kj���l����v����ӗj�k�w� r�|C ��:-|V�h��m���O�G��B��cw���Ӿ��Фhf����u��m��m�E����.��������f� .����e�^҇����fC�P��"=hp�"�����Ҁ�"d�� cge����F,n뱟:e��yy�"��w�gz%$魼�� h⊹��#����Bl�N��%N�XoG���w���ȑ���L������\tV�r�Ǳ���뚝����zQ�mgJ�dH7�,G��oc�'�O'M�hl�j4jA�W�T���������p�԰�d�������w������k��>5$���\z�f���۬ǡ�ǧ�曢Od��MDA��FɱM�	6b�>zH�Į������'.{����a����\ �h�ς'����ː�5����o��!I;csѥDd 
��ܘkJo�N��f��J�\&���,;:}x��k�@9���˭��Z�؃���b���#Q��~لc���#�Ã"�f�v����HG�aT1 ��=�mqgf�k��-���J-�����Ň� �L䈢��=������A�5�a���@��5z$#��)�V��!dʸ������M�'���΍���(���� ���]�-�	������X�'�'��Z��f`���`2s�B#(pa�x2����ms�b��a�B1c#R��F�EiY �����fa�(B����l��_k�u���%qJz�j�acLR�̘�6dWa|C�rV���Z1�Qvl�D���q\�e���ю�rf���a�>��l�瀳
�a�$�ҧ{j�i����%+��ámĜ k��.�aZѥ����G)���%C卾��{���%�*�)7�^�Ź�y��yjc���Ӣ�W�������S)��V�'[�������Đ�o�1�@T�m�S�A��cy��;�7������	G�dZ��D���]'�.��.l���r��t҉��c^*����3��9��Z$%�$q���d@�Ì��'$M��Hy�ԙ��.bGR��cµ�⩼�)��a/����0s&�St����EK���8���v� !��,{�>�j@�b��D��������12J֐!�E�$�r�
-�lnɮ�� 	����#e�����HQ�A�yDqŹ��m�������n������)����������K��o�wE�0dy��L��Iӂ�����$z"A�B �������@��Q����`�'���uT��
�B��%m�`���X�%����:gT��e���tí{���ȴ�s�u�D8]��d�%���~������������me�V������S���}R���h�ʹ2�9��Ԓ��T8ԑ�ʩK��s%6�wo