I�^�l�����xe��@���c���8E�9B�>C�?D�8E�_�{��W�..�۵L1Zd�O�럷�w�p��'lхaĻUJ�Ab���ڜ���Р �0Uߺt�&?}�Ԉ����ŋ�F,S��?��g���q��%]T�"GNJ�rգYα��B��K_>t�x�P)&�M��	!�`��p�=@7�8����ͧ�t_?�OK3d/G���2no��|w!@Z��\`���45Y��8Ta��)ͅ8�Y���l�J��tyC��f��}b�-q-w��[c*���ӻ]���ȷ;��R���r�+�=vʘ|-���:�<�h���p��ޭ�?!bkhf)khy	k��T�~�V�~Һ�,%�c%��\�[��b�[+����,��?�=`n{Xu`���= �)�V���*�`�t��ek/��J���Na�O f�B���<i��B��/~٘/~0�b
"��5�O-@�~_���K��QLM���S8*�����L3���8�zgA�,��|s'P驄�fG�@�l!&j�Ŝ!��OH�7�����yk��i����6C	+�L��������>l�`U��.�Ix|C���@�"_���.�ʍ��[޻�����r��z����n�_ä��o�j�=�ΝV�.y��dgD
���ey��Vel^��ɖ�Gh"'��M�\
u������Z4��<�Q�\��lDZ���SP%}�|�d%\��|MY+�1��O�ѱ��]���I�׷�����ov�xdc��k�����f�pd��"��ס��)��3�\���^�����O��曶�w�
auN����3�gL��!�쒹-�B_�9���}ڱ����wi�k����Yf�"��'�D	�grK�U�P����K���}�n~��Sa���%��nEǵ`Ŷ�}e~գ�TLnh�Sˍ���D$,��Gt�|���%�|1/QȏS���K0��r�ט��z�,�wT�s���y�j���of �]K�`��7U���NZ�A�s2Ϩ�v7���x:|��0j���"��FI�7~�R�)��t=b[3�ZS�1�Ȉԉ���Ϣ0���!W>�����m���䜂k�J���> �;���a3_`�<����R�Jr��=�2�%v 'ଊO�-�ؘ<�$�4�9!檬�TZP��[|��}�;~�f;|�~;�<*��	�l�\��ۖZ��K�5u)��C0�Jh��
-s[IB��	��H:p\AeM0//�Z��y3��|�F})F����Ժ�U��S���"�
��q��i��/��T�l� F聆LC�O��!�h����]�!Yl���k����z1rԭmժlҫ��ݫ��E#�4��5��f#� �é7���ǵ��)�ҰST��t&�4�(���?s�,�π��ȦX���ql������B� %,{��HWP�`��m�1q�&�䱯Qo���M	��Ϭ�q�?k��@Υ�Ve׍uYJv�F</��Y!�J9�,��={��D��`C6���:��uVV��h&ė���kؼ��04;�o���4�<�D��[�#���e�\b� w�f����_4����|̉%����������Z"Z�3Y"���[$�s���@!� ��A�P�큻��&Ms$��
�bb֓�79��xm����,\C��^�jዉz÷��x>���2H��>E��~�9[ue_)�j�i������7B�Sh����Y�9��r�7z���b�[cS�e�]oD*����1*-dʥ�
k�g5�>����sJ�s�i��3��۸ƿ�E0M�G&Ok8y�Z���u�x� 
|�����d)4���K�&���`?�y����s�ӡwaA��q*^4{�jx�0ӿ
�g�V����J}%���]���`�èZ�wR������1�r��hK�r�H����>�	��w��E��2�����ß�����f|�#	%���ʮ������r��cE��駄��b-���~����!%T���8��$%T�+�0k+�#|D�\"��b4��z�)�-��TǤ�\��nO��dx|�R�#��(Qe�~� ��ؔ

�Ք$��\�	m�mI���>T._���.���@:���d�����0��ƛL�t��#?A��!�d�"H���'����iJ�T�a�::�f���7�+/�k���5c�Ti�eȦPE�9�z�������M��)����0����Ίr<1��:L�_W�Xp5�%+��G�'o�=(m�*�J��:O�)~ɤ��z<��*������u��P0~�vځ4nN���W����*����@П�31�4���(y�E҆]�:]��.��Fsf���lK���K�ht��sb�d/6k��ዙ#{�$�o넘$z��<�����灣 ͎6�#�Z��<��?�a����p"��^_mdu���Ơ(�9��d�x����r��`����je�5�0n�l�����u�$T���14;�|@�?U�Y�uY��҃`���n�]0Ê�A�s��o#	���=V�Mx��/s��{(���n$��Z����h�5;a���ba��ba�U���괙C##Y�=~�Ԣr^͕�Y}s=���F�p��Ik*�"�F;)|Zq���lY_򉱾��A5Zy����c�#����T��� RX���?md�0qyF�x�4�Z��s�8�ș�ã,c&�(��~��=�%Db���ځT"�Fp���@�j_q�Z�����.����ņ%6�u��z�t�'℔�d�������d!р������#Xt�����P��0LrI�R8�fN2މ~�����!�]t�w�%���`u���kƫ���h"Ȭ�[����RP��ٹ��H�#�Τ�����n�ܽ��?�Ƀ��2g8�����琊wh����kr�}?�u�u1�|�ae�'j*r��ѫ��z���o���e	"�5�d��<�k3ۜ��8����nܚ�#������c����*��Cۛ�"�u��DE�+$��ʋm�c�ue#PA��0���2�r������@��}���,��š��~�~]x� Z�������2�a� CU��A���A������5�g�%�A�d#���]_��Tr�����x"Ϭ[��}��t�m%��:/�^�n����hm��[�Qs⫵市����W7Se3`g%�s����X�[
�_Vy#��4��r�Ѣ?St�C��a���O&�[s�eF���$�S�����o����H����Ba�9d��zP���q�U;���l���M�¢܆��f�n`��<i]�,��=��¯�����b���eX�=�m�T>0�u��=�cйIs�cI1�֠/.b����?8���.;ܴ��J2!�����?�點�?�Ef?��
�c����q,X�&�HT�`�R�5�����Na
C��W�#u?��� 
�hϳ���c�9�K��n�dz�*{��+7��-���HS��{(�
���P�X��6Ju������.�o��
۾��;�Ӊ\���[���\����[~��x��(���+)� Hmbq"p����zV�q�F,�����Z�bm9�%�;�Z��A<n��tQ�4ѐ�p�Yh�,'���U��.�4�������&yz�Z��i/�������1{�M��Qw�e���t����0�����2=Ħ�櫝����.�c�������g����ٛ��Be&{�X�׹�6'�s�n\��Р�g������c������n]�+Xa���{�דz漖yԡ�-�1;o�c�˞��@%kB�DnJ�ڵ����)��]��RZ}�y�a�D8K#ܱ�u��О�6�?xNlnhxiy��P�eb�H�4
yn���6��y���K=E����1��1�J$��v�|Sa�������Q��7P'�t"6��0��cѰ�K�aW��U�nØ.�<�5!w���|=���u��dli^�pI���϶�V�::|)��A�Q��;�7��Ku�N_(�([��������3m(:��Fc2���^��E ��Zn�~8CI�K�FŇ�r�X��^1��T�4��|V���As>J������8�����8������o1�}ĳ�ɨ*~M��.TǯBm�����(�^X�;�,��O%X\^�25Xs���i�\w��(�h͏o�9�5Ȍ����E��@�|/Ip���Ak�pw�XN�;���0�H
h�*-�R;M�6i}���>�3S��ñ
ʷ��]D���ih!�V���y��3��#��vU�H��)��'���nq�/HqZA�c�1��kI6�M@�&D:��νF�>�q\�o�M�����)F�N�E8��ՠ�IlDru�U��wQ�.$`�*�Z����H��P J�h��xw��-P����%쬔a~9*�p�f� �Ȋ-P�,W�+V�*Q�-P����|�4���\m[
�NUt��ׁg2�&���J�|F..7Gm]�"�1l�2����՛B�'*�k��P �Fa��Zh�&��SWte�����l����9j[�i��J1��
]�#�Ub��>��3����3�]b����:�^g��T����`1V1ҭ�3ȩ�Γ�'tkމi����9=��^8MU���"q2�#{n�H6a/y��F0*=�D��'N�W�j̺�T���1Rn睿9O����Zȷ�W!1�q�f�D�qnǧ;���������;2������^$�"s����# :�_�	�(��g���tC�p<��ފĩv>*�CV�h�g-JF\Ξע�H��ʀ���(h)Ѡ���]<:x���Z5�	N]��2��TnЛl[;�i��o��!���&�8�B����ȧ�far���nc#'�c�6�f4�02�' w#�/pPvd�����G�ĵ�ϧS�И�:�"`��I��l7_����Ɲ���_���!���a���#)Z��g�k
e�
 ��������U������R��g5�>M�Sxn�)P�RD�����j	ʮ)��K��!����1cs&Ĩ�/Z��gi1_�N���Z�F����Z��'�_9|��V�ڲ��yNt�z�I����h�K	JXd��K۵�UU�7<о�p�z���3��;��,X~ص��H#]�� }Mt��ߓ�=����i��b�|�lΗ��kY>�
��G�g;����t��=�-����O��1��Jln7�z,�e���p�!Pں��F����X�J��v�'d�H>�ża�&X�{�g���9_�g�橷� ���;��������w�:�1��-���?X��p�xe�)s�o�x����63��Ikd�m�g�/U�b%�O����V���/�DAO��F������ ��_&j�ǧ��mX񠂩�z���Cg���8`�4>��Ķ��71T���?{������A|CZ%������Љ�Z�ߵRѺ@	��<Z��8�ɒS����hG���Z3��m��h���樠�4�T�蘸��2@H�@%	��f�*,"���ĉ�}�s^��͚������<a��;��`��،\�O��lO뛠}b䞂rm�42�<u�	�Ȑ�|����rK�P���غ�pwO��j>�8-e��<�k��z��.mh]���.����]"�K��w�K��x�Q�p,�����|���ty[]0�����F�D�s�F��q�ɂ��c]�=����ZO�a�(�H^J&{J&�\�aRQH&�zaEӟ��E�b1��8�c��Q-l��\'������n���ΰ�O��zP��.��\8��^�ݹ�	˼YǬ������S���� ��l����ťu�m��!
�9���E��p�AfZ���&uM�f��ӟ�h�Hv��6�(ꄆ��#�d蘦��L�Ku��YE"U|������]0o)���?�k���� ���}-F�sM�mm���r�%���6j�f��pD!��O^"hl��"� ���aJ�gRI��C*gg���Ypb`�#��Ha'�q�}� �Z8�/�^��2C'