��������������������$$������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������ff����vv��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������@@��..��..��..��,,����  ��99����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������,,������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ����    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ���    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ��� ���    �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���� ��� ��� ��� ��� ���    �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ���� ��� ��� ���         TRUEVISION-XFILE.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                < K  ��� ��� ��� ���    �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ���� ��� ��� ��� ��� ���    �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���� ��� ���    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ���    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ����    �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@@������++����������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""������!!����������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������xx��  ��ll��������������

��@@��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;;��  ����������������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������qq��  ��@@����������QQ����@@��������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������44����**��44��

��%%������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%%��..����������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������cc��  ��JJ����������������$$��������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������11��  ����������������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������88��  ����������������������������������   �   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������xx��  ��44����������[[����DD��������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������&&��  ������  ��������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ll��bb��ff��ee����������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  