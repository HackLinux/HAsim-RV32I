A(u>(ׄN�6�o�X�f��7�j$ �[�D/��\��#���7W�i����.YA�UkJ͟i
�@��Ғ+Ճr�l��\�|m����'�6ù?�����o�(�:X.8׽�y`2	�|�.e���(T�}٫�6wE+ޠ�j��||.8��n�@��7*�i#�XZR�>��C��A�x�y����~�\�� �u)�����s*���ߠ�'�N��Kb��%dsXvr�i�
rw^�K�a���2��z��/x�S����/K��n�?(3�&i~%T�+i�Ǿ�kx*⡸Nc�AoV�����k�n�����H�,�Ҫ{r��&�W�n�$+�����ej^O�Fk�J��_ j�n2w��J�o�6��3fL޵H9�~����|E�X�I �y-���\�V�(��}�����V��)~�\b
j���^��x�k��&��>��(��6��a�j3���dl��c�Eo�l#-�FE���,��j&�G})՜���[rr#wR&��-\�B�Ք�n���(����Z�&{>�ėd%~a��Z@	�/k���D��EV�E"ϭPW�[�1<{�ϑ��,C���*4���y��|������T����j�9~�b��x�U�>-%�+Bs˻'C�߮��N��aИ
�L�u=��=7���1-��1ȵ�'���������PZs\���<��ߘm����4ީ���$���q�Dz�NҤ ,Di����@��/$�ᘨ��%�j(��$c�ם�Qs'*��0yx��=�&%Ġd��T�/�̌��x��	���2�!_Á��F�u��'5��n��ߪG���T`ۤ�FT�Ӏ��M���b��O>��.n�`l$ӥ�j��閣�ڀ���X)��"*���T��h�F��2̛�C��ŭỴ���&&4�,�T�nu
�{�P��Y��다AvE�,��+���)D��B��k1��S�E,p(f�УD��|e�������*$�qQ�3����5���إf�֑	�����R��
�(is�A�:6H�椞gꊬm:Zr�r$L�f�@���2����]M4��G劻� '�)l2_�ǿ�׌�j�B3�9��b�����*��$w��aUwr��Ժ�V#Gg*���*!Y��VR%�C�>i^S���9�1�Ɏ� R%�m����3?�W9V�L�ē{���0�5n>/��u4V׆Ae���ȺUl�kbx.?��=%�Ya��<yi��8S�&�a�A���e���;�����z��6���;�����&"҆`�<-���98�ov��,��h�bHhUa�aEK��$2��O �G�sx�	�1��K������_2�
¬�y�SQ.Z��P^M�/����ǂf��)
��!�q9�N����|�����}j�3���}R!����¢�:!h�����l�8�q�<���/��u�Xr`֋*���\��i���n��������h�'��~�9�0~��BE|�J��x�f��K�H�jd�l�5��e�9eW�te�cd�)K5�O9�4���?���h��8J�sP��u�~�z�3��8���-�����)ڌ�u��Ƶ*'�e�A�6�|3TZ�k\�R�r�m��ÆB-䴘��0\�18=��ґ�F��+�GA����h�1�峿i��������+�	mc�	*�_)���(�,��"�Т�e3��/Wc��oft&���v��E�A��!U��	r�(P�G&�!��Z�'jCWc���-�-�Wo6���+}GC��U�J���V���e��r����5�L1#�Z���� ,w�鯍�A�ڣ[�)GT]r�98%�ՋS�����.g�*�mc��C��3A�L���)��[�K�3�d`'5����	ޒ �L��8g�e]K�Ҹ���bl��}��Y�b$f��MOB�\D�0��(��3�h����9�͌����r"�!��ev���]z��\7�#�U�爫u�N�XS-xa0e@�
�ܑ�Č��[������6����q����G>w��cf�k<�Ջ(��i1����P�}g�fE������P��:V� ����꩛���� p
���3�E�3~�J��{-Y���ͫ8��V�T�(>q��E�k��F܈Q�&U�>y�D�0��AW��@w�)3|�jb��Ut7�rKn)����)���(g�<ʭ�X�ˏk�8T=�+Ѿjz��1d�����8}1d�愺�V�Z�bq�z�i��&C�����iQ�������R�d��c���0�ҀtԈE����?K�/�����G����z�繸D�L�������i�~-�=�B�lRp���7Iһ�D�P�'Y�� ;���Z`�7�o�(
�ꎻW�/ޛ��l6 Ux��c�:���Dt��U-����g���߃�bX2� D�:vN����qŝd�����p�b��-X��?*�"9wã��)��L�D�f�e��W��ΪB��������-��B��"=�a�24~���a�����5�Q�q�(eD��7,6��~�꺠t䤄;��:�[����s5�>��Eya�D�A"~q�_,���`��`���rQo*��>ac� :|��ö������_�'fPwi|G��WzS#�U������ڎ�qj�����X����ۺ��c>_q�m��U�@��6���~b�l���=������t�jE4/��|���7�V�xmK���p�T����g�N����j��A����FHr͎lE��x�,��7�"�N�	���.���Yǒ��,�#�w�]0�ĭ�$Y�z�R��+�.0$���~o$3N��ԡ��t�uۏ�b3~���@.�q�wY@��9"M��9�0�(B��`~^����6�����ɢ�k�,"�D�a�w�眷��f^Rݻ�s�f?撬8��Ǹ�z�����n	���hZ��ϴv�t����������Z����JV�̏��4Ye,J<>�
G�������X� ����4ࠆ�G�t�:��Sx�f=�7�n4j��$�2.z���D������^�1;!a{��x�k���e�瑤��q�*���q�����qϐ�����Bɞ͏�y���sRuj��Z\��SG�;�-RU�ie�.�N�Ƒc󐬝�M�T����sq�v@x{Ǣ�r+�5�#c�9�*��Q�K{h�����r�h��"��a�������~����Ŗ$�]�LIO4���"��}���Ρ=d�ВbpB4e[;MG���$뗼���؋n2{����~vR�o��ٟPáP�љn����:߂��m��<�k��1,�)�E�-�)L���s.Ʃs�E������m��HB��J:b��p���ǧ�`>�~�h@�n�?�������Ť"Mƽ��kk�j�2�.y\GG�~�+�x�:���t��ޤ�������Z �Y �A�܋�M�t���sm?�rwG�������9M�IE$��6�(�^t���I��Zjm������,�f��/B��`���w)5��3�L?�T�&���5;�mL-�����"�C�_�'�Q�6\�d+�ˮ�%�G�VEB�T��쮑�@*FF0���o*�ܕ�&V�ň*����H%d���R�$@�1ր���VQj-����r��LZ���uQ����9R�D���`6���maf-����B�a[F^`�4S4���Y&Rb$BY�x� V7ؘ����2X����� )�G���unWy���t��oB-z�/��l.g��2�������kC�B�xd�h���[y4��ɑ�����Sz�0�4cod�d��c�d��E%������B��~yVF�'���EϡS"B�-���0�}��������l�lD��ĪFF��M���4�����֩�ی�"���x�!4�5�:��fg�� ��'$�2���4���Ҏ�gp7e�x��|�G-���ٻl���o��� TnD��n�FP�j"W^�ݫ-Eq�B���� g��"�}s3}|t�~��{�i�B�+$���E/��X������&x�Y�e�������7
�ndWZW�+2�U����my�=����D9]�m�g9�[��ڔ�mcp����� L�d���q|_[����>�oX7�U88�E��n����/��c��U;`�@4��	C�a���Ϡ��1��Q����eV�j�t��9�'s'���,��������R��u��t��)5r�*��(�_|('+z�at�`sO㐩�<F:B�2�if�0��������L�.ٹ��~��ԗ~�ya f��`�I�&"�ϝ6Z��3����d�vD���P��W�O�U.rU������u��]g3�f4�"��ƃ�7�l���l JĐ4���Rㅳ퇫a���h4�i���͇�7�K����X�4���3�	�S��)�'�N��I��\�+�r�G�@Ӽ��{LO�dL/L���~Љ�W��xă]Å����@�F��`�N{��5.L�9��	���!�V�2PþQzX�{�}3�����6H�m��_7pV� �X�O��H��յ-�U9r0�@���[7/8����^����,�o������3�4��*R��j�#r����d/�P��/�Q���Mn�c��dw(��Fp~��\JF���:�k*x"@}����� �3X0{H/�7Q�C�<4��&���?�ਝ�i_61I���M�z�/�ե��C�@�o�����Uᦏ�jU�%U��Gg�RyMV�H1���D�$�9q�l�6TP�.�5�+��X�$@U����=���!��J�Μ�爫ծƃ�r}cTh��#�X�X5��k��j�ڏ̜�e'C�z��n�i�ٵ_��S�f(AP��vpUq
����RK[�<��QL�/%}�@�Y���_!�+���Eި�����^�����I��H֦��N	��"A�l<�X�	��g<��r�3L���c��v��,	�����\.AůߋUZ@ ��	�%��"�y��Y!�M������))�cT�����v��B��v2E#��:E7t�Mv{Q�>�L��8%@��lj;����;+���3CٙD��LyAl��ՠB���[�]̈́��[��,���]p� ��ҜO���vJ@�#��!MY3�<`<��z9MKJ�a0�����L�&�%�����Yj`2�"f|?Lk����D���v}���层�ETb�6��T�f3��kG��#���[��zo{w�-,Hu��Мd�Y�sӇ��s�/�kQ�D�j�Qn*���^&!L��� o�P�E׽k��:���Q���.��/���K�炬rǪ���|"��-��|��C���e�94̊�kdX'���0/�[�Zw���	��N��[��=�,8�����Q�����m������j�~`�Da���<&�E)�;�����b� ݠkF��e`[baL�d�J�wU�2ea�'�Z'�H�����b��p�>�G~�-���B�!�no�i-��ۉ��Y{�~���!�\x�a]#f|�b�(��,6�l5�m��k��0i)������hW��.^�~ *�ú­4�l��V�]�~y�i~�-\>Y
�K�&P)H�!s�-4<O3=pz06O:��\�{j�'���0D��a��Q�1��u�5����N
.����Wc{� �+�j����C�7�Ψ's�(�@�����i��3�Ư�ǨY{�o�����Kj�ֳBH�iUz�x�i��j�A;�3�"~��t+�z+d�(c��v�UDc���J�D�-A�M^��]��Z���?��@�cx`#xa�i���& $������������������*���"�@OÖ ��/�&-<4?4΁�Nl���5�~�K�������K5���щ����w���Xf���HUwP�`J9m�'|X�����i\CEz٨��=�G���?�	��L'�^�Vᴽ೬�꼚�A8O���� bמ��ܝ@W�G����R7��R�!�ΪX���æ�Z��}"a����,]��_g�gqc�4��G� ,�ߪ�8��A������U�r��Q�0M
-\V��8�Voyd\���5x�i�7����ݠ���{��)��(��{<���3چf/�k���9���`���B���/��h�;0�J<N;=�<��b���"��%�9L�i*�H�~�o��
��oh�.�I�f|F�2�_��UC��