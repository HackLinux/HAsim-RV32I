ߣ��ek�*kt�{z��[�r�6�g����л�9�Č��WTlyxx,�YF��n��;n�[���lM朖�\c,��[Xn:7�Q���������l�[oxN�a|�w���,����ϻ��c�J�'l����Tq5w<�a�K�I�QJ��:��8w�{l6�6�~��T�O[(z>/�H���7�o�848_�F�-3��P��F�ҳf��3#s�������C7R>��r-�SEkf��~���=s�<5S6I��+gb�\њ�o��!�X�ZnVD%d���AP�`�ݙ���1���5*��8���26�q@��,�&OX��,vH<�!ۙ!e~F�*6�h�H��!bb�8���E 4���bk��
E�~.��(N<�i�Eϥ}���CX���	-P)���qB��棯 8�t�u�ȸ�f;����Er��y�����&7��#�]��~�ʟ��<�9�K��I��&>���c���z=�y�pV�<_S^�#�A�Yk$���x�͢A	��h��ѾS��͸ ��XC*�S2Vw�%��G�0����WۥW!g����V��W��}x=���xl�]�������Ϳ�lh�A��S(��-l4Fwv�����ɏ�bA�˞Y+�k�e�nRGO�_y�z���Л�1�h��H�,|`yBցw3�D<�C23�Tk	5)�[�x�<x�z�X4����x��8i�	����v�T�����譠���wq�Pj.u� �Vay�Lb՗���l'��3)���vkg���6�Y�aG�v�f��h��Y���42�׻�l���uя��[씽��:֯>��p?�3�>3� "��]0ؔuRX��Ҡ�C惦8O.�E��C�lV�!ea�����*��w��3)�J���\��ּs�ϫ^܁�ѷj�A>�8'Yݑ"����3a�\c�,e�_~o6w9c�fA^/�;��^G~W���XԆy��m��oW۪b8��|�r$��V1��!�fE�3h�K�)�Qm��VFN`CQ"�%��w`G 9d�O�8ۃ1{�P	I������.��{���ݘ��h��]L>���6�z�4��-���RY����`��X���i��^�%}�K��A��åz�ӟ�����C�ϟ��&t+^Q��QL;c1s��[a�>���]����(t%���O����ߘ$��H����K�N�0a#�Q���������|���ϤP��߶8�u��+�i�ƽ��C:7-O��b�ETj��z8�~1��-���V�L�{ŀ{����5� mM��$�A���~)!o=#��Y?lŻ�-��ӻ�˚<C���mOTno>��H����/��5�����5�rz�����U|r%|/FA_.|6mv.�9"I6״+T�Ѐ�\j�a�ұ�}����O�.\�^Q��7��wh��G�|#���6n�}<�2q�R���G(��_��mo��y��#Cص���´����LpN/���x3�}&�l@�n_�G y���zEG�z�[��혰�"$�Ζ<���6$z�x��?�w��u�Bo�H�
>��;.�u�{I���Ku�� m��l��Vd>�9�]+�G�U[�M��!h��sn���;C5�܅:�1�:]��U�����*�=Gm�i$��}�����*�l*��S31�c�z��9@���kc�1�zQ}LR���nU7��eZ���� ��V�u[�<l�{\�;�E,�p���ا� ��h�iD��Gc|S��n$�%a�G���"ֱ�pc`�!6n��̸D��63nz7R����8V�z�2���&��b���,>�, �6jYfɺ6�a��hJ֦(���+����W��08vJ��u
bXmD���ul
GE\��0�	As��|�1��5aV6���Zhtͨ镲y�h��d8WHZdl{A_G�ӗ�
�~��p����$�A!���(m�8r!o�y ����L�9��f:�l��B�.9N}��>5䋱6SXA��T�d_Y;++�x��C_$"1�0x�,m��:�LL�����}�/#���pc����.��2K��y#�����\Y�+�q/�2z����oR؈��\a����-�y�u�����/9��@g�
놆��+�6&ê��к��%7�$�pZ�	"8% ���Gt��T����"z��>�̠V��յ�3�?%�6;�7j���rw��I)h�����-�	�K�]gÿ�G�qg0j�z`\��r2!2Ig��/�N�����X�+c�&�5��+��?��7��ț%:���Y��~�H�)X׀_�P�ݧ�\�b��5oL���i�W��8мm3��yy?2��y0}ޙ�/�ug�^���-+���&;~������#^qQ��},��7��a�����4V�l��'7�i�|٫q��QD���i��j�Q��$Gm��V�/y�s1����۷y�F�_s��-�z���H���?�{fx޷B&��DN\d�K��߱�Yds�}���-�Rـ4Ԣ���ӄ�H8�B	� ���t�q *����+����%7��Wg-�rjJ��&s��(�G����d��w�u�n�}9��m�9���ʬ��>~�Z�=��l>�.�
�q�(�l�j�#z�Y4�fe���̀�nI��8�K!sɋ;M�A񙾀�,Y_�@�w@�����$���+�@�ei�`6&�
e���T�Ixi���aK���rC 'ѻ��m[�)��Ǫ�h�ۊu�&P�ُz��C��,�m��6C�}V?��<��	�S3�2��+�����>���Y��	U��L���.��mQ�+ _M��&��Eia�Z�ET^b�`�{�k["�S�U;�\P���$ۑ�}���#�������T�BJ̮��U}Zi�CEH�e)����aV�[��X��f���N��.@6H��^���7�ؗa�j�f�Pn�x'���2oTV����TT��x,x��O5F���hw �d.7�m{�z�� Z"��W����1$��Ύ�����D�B͔d�2��@�uO�����=z㴷����xܑ_��!zPt��q���žpu�9����~H��N&�9ƽI��'i`U�� �
\�*�Q릇L[��d��ӥz�n�Բ�.�\~<{ǹX|��55-���%���e�Ě{��o�?:�����J�
πwXFƠ]f2�#�_18w���pLR��8L��(�P9�+�;0|��'K%C9AZ�y9�#6I��&����J��3���Y���B���҈��t��5ϙ�Hb�u2�9���5���'�Gvۭ�����!�a�@�x��$���ت\��:`����̞v���՗�Q�شx�h[w�`$@Q��7E읱O���O�-#R���԰4d>�E���{�/��P�%_N@��m��U�X�$S,j�a�B��jF7��c1�밙hpۿ�	�	���
�5PeBu����4�+5��뻹60f���VˣRQ�Zdx��TO�|�ޠ5Hr�\N�?2�SOD�[.�{T�/�aH>��i� `Ҵ]k�Jg�����eù]��5�M�H�B�,R1�w����d�����1n*�,�YV1�H��"�ݓe�?1�9/�WA�>�j�r���-���_E����IJm8S/i�@���X��e�M?#L� Z��v)�e�Y�$%V��o��:�\��ȋxe��9l4|�$�����7� ��ڻ��dg�C�ju֎jM\%e͉j��V0�Q�?i6_�i�F�y�M��|ݑj/��|ɵ���^s����\c��@�e�H��)<��慴v���f��z��Ǫ@C���0D���|?���r�Z�Q�Y���8DZ��D]6���cd�g��K+��������Lz���R��Z:�g�mu)��q���L%�dTR8�Nhu^d$�-���|{�|�|���yh�)H?�$�|�������!�1� N29Y��2����ԃe�8mq��/n�M��ͅ嗣\�jNq����M:NJ�uU�&��b��D!Ț��j��G%��[�ꢖ�ߪ%�Ǧ�tC�G5�?�.u�������J�^ᘺ�>5�?�&���[h71y��b���'%S��Y��fl,��Z`/,�IoE�e0�=�h��xzD@���2�u*"+U��l��O%S�j)��j���:io�\�"m-�*��ʍ��ʬ�ׇ����x	|?́P���--,�ź)#��B��xWE�Md�=�U1�y8����5id8�.B�k�</�Τ8R��ut���/��6�yʡ��� �� ����������������WE�zܠ�&�!��/�_�����A�ڠH��� V�ߌ˧�� E�d�;��K~6H�rjPT����1p�X�z���3����TmSr�f�l�Sн��jLKM�@����e���Ze����HP��(�F�w7N I-��a��v2�ui)����v�
����n�f�X�l#�YǍ>�w&'�|��C���Q7���%�b	�gn?�|�.�l�RZ���\��sR1�]�(���\�i��E�bY`��@��a��+��X|�M�چF���zN�V2S�	ra8G(s�C�c��VUt~f_�(��5N&d���Т��c`rD�w�9v�7[�py��7���UI�ǐ�¡�p��۷T���mz|��F��z���U;.ϖ�|�����$`��.X$�{'�j����rJ&م�uiV����,�s*�� (��9A*�Rѥ��R)׹D�թ�<�,��$@��#�.�S��|��e_'ғ��L�w)ɥ�����,"�]�QL) /���d���~��i���/���c�5���x����}����Z��L@��8�ӷ�4��Q�r�7�261ҍ�5�Ws'�[��Υ8E�T�D4�Ƃ�-	��"���J�jPwRaKeQ�����W�YcC�"��/��ȓ� �$�*�@�Te���50-�ɘ3+8����	r,0�!2�J�](<ouɂ�Sќ��䟓� S:KJ�'�!:�5�=B�Bc�u����Q|x�˼��2�]I��Q��P�VJ<Eߩ�P��	��ӟBD�eA���l��0?
Vy������q<��SVPz���֋�'_�����F�dD� �(�oҌ�"�K�a��y�����5ŎZ���=��?���{��LR$��2�Obe�dwٛ�����ؽ���V�n���F�6����ă<>Lډ��=������� j���N�0:����9�[���d��ϔ�`AX�}�/����ޗX�1��;�, ��pAf�ؤ������y�� �	6��aG0x�m�>�K\Bhn�h�C�����o3�ą�O���WD�-�D%F�~�x�$�ޔ�g��m�V�xC��o
Low�x8UPp�p��n��@����!�XY�,�G0��r��~�0#�^��M����W?��,�g���_�0ZuU��=�/v&�WH�8k<ʘ������D[��?O��(7�s�/�I"1_/۶>�08��l|<�P���~81��D�|q�bQ��`~�w��p�A��Mg���L�<\�x)t&���76����qT�`����9�G/��A��vT"�*?�ԯ� ��1w��EĉN!dg(W�l?��l�pl3²��$�b�!�k��yW6���(�KU$�D����I�)�.���~v��X1��&Ef~g2�2ە�/)vI~�3nn.kK�c�\����,�I~ŔS�,m+��p���LeH�F�C��Z0�� 3|������=_�����?J��� \�~.�y&�s�s��M�Y�7�0�z5�Qr��M+����IZ~*��=�xl�ɜ�����!iUa���|�Y���w�Z��!Z�z��PbLW�Ə�p�j��Y�i"���/�Ֆ于��g�@�D꽞��$�$N�D�35?��O�L� t-�=xF���gՙ�@�����D5��j�T��g��,�{Ѿ_��q yY�{EL+!r�g�!��=d��I���ϓr�����߅O��T;A?����q�!�|�]!rZ#��:M4
=��f��'����
1���<`9�]��f,�<��S2mN~l���g���uuL�o��f_����%���e���ȗ�iFK_�C�,�}�Z��]�:4����l��n��i_3Ʃ��g�'��������^錴���)1�	�+�:���NG�����<������v��ǖ�#w=�9�w�e�ջl*
j6������f�M����<�����^ �5{
;�;��$���VC�bR�|$g�ڼe<ä�s������p9(��_���9�c�Հ��x�N#p�=i~�E*K���(���Q�x&s!,IW��荏�Y@J#�
��)m9����,cH~�P�����y]�:�jO�,�$V�zÔ��T�|������4}���1󳞴3C�6}j]Z7�-��*S�`�Ի;���@:d>GSi#�N�;�"��j�r)�:�f*W�3��Ɏ��Xq=ط�%�,�.95�{�ۊ#��7繾��eu�>��)w,�40��TB������F�ҾFNW�5G�V���z��K����'\b9q<� ���T\��m�����kZŝ�F�5%�������ֲo��uu�ث��u�]���nu&/�c���4����=�@n�H�i_�T�Q[��V�9=Aq��6�I�M�+=\����v��h�\@lg�%�u���W�	B�Ʌ墻�e��יW���.~����5������>�E�W7%ʌ��?��^��a$�F�I�w�>�\��\�Y���Fq�T�k�1Yb������d�C��A��c�s��Y�ahz�����y���x�v	����$:�B�Y\��u��-����g(j'��.J�a����u��I�*ȕn�!����Nuu�a��7K��H�N��F�̬�Di|�-��9��u���X�ܲ�O�m�`j�hZ�l�����>-���OG�U�m�^��Tp�ahr�G����J����[̧~��_R����r�r�S��ɘ�`�	W(�Gkf?�tȊ�ϣ,nno���4ꃜ�&U��`���V�����(�>�82�ĸ���g$����хY�0��>J�ϼ@��~;�;o�#�g����ѹ���D�8_����=�z]��q��i��
���}��H�0��B�Bi�yꥈ�ZO[?�;v��t���?v�P�\�~���8{�L'�y�ۢv���s.���,Y��
�Z���[��?�yq'�Rr;�5���o�H��,�(S��j��`<�8.0�[�^|˳h
ic'Z�l�͜Wpe+�	�n�����H�V,�J;���qB�m	ʽ��ŬNl�ϭf�+\<n!7�~��������S��.����U(�c���=]�ԧt�x,Um�Nm�,����y�x*��K�s5����<�-����{ŕ��=�|�y
Hheg=���'F��fu����Q�2��C���]�
Y�Df�7�'ɏ� r��D0@Orm���K8�F����D{��ɲ�M箧��#�@�EN�9s�i��W���&-�=ob�֏��\&ZԬx[��r�~��o���8���M>D�چ�3��E#��M��f��� 1ɞwV�N���̯Y@��%{�6�M�5F���r�# `����RAu;��!��S�&E�Ž=w���=*��%��I,�������0�f�glO��u2M�\�����N�Fzl�����]* �U�a�D��-�/Ɠ���Y��E�Q�����[!Yn72�==g�(�҈�B4�����U���St|��CJƀv4$�ý¥b�Y�
��;��-��ַ<�j^���?�T,�^[]�U�FLh:.�����ti ��G"�)����)8�G�
,��
d�W��t��8Ӗ|�h<V)ųkf��!k��+P?�X�"G���|'v�A��*Y>�2?U��U�����X���������wҐ�\�������3g|ٚm'�I��[mO�����|n�G�zi0K��Hv�V��ϻj����nm�vn����F�˹��i�}D	|�f�|�[�x�ʙﺜύ����S��l�>�4O���N�8�=I
�I���'�LFo��G������I�
����{4���א��6y�����OX|2>�hH�&Ѯ�ޣy�A�����ڣ��h�Qƪ ���b�L��D�z�n��E^��"�����h㑬;4�GE�'���r��mMf�a$��4]�r��?L+v`��P�jQ����P[*wN��:s��d�bP��h��]o��(��۰2�f+>�qc��Π*N��F����V�ξg��@`�@���f�ɯ��x�1�\�n1�.��ML�gĢ�}w/	�,�u�����1r״UC�k/K�H�2^3V=���aXS�!f9��a}lغ��=��݇�(��� ����K���.���\1����G/�ţB�{cz����*l0>��E����]p��0(X��5eu���y \a� 8���7�f�=ID[8-���W���$��KԱP�5+����������ݫ�T��0�����h��2�My\s��DkyoL��[�HR6!+(�t�ǉ�z��̼$C
6�I� X�.�z� ��<��ծBkM|��,䣠�r�B�)[�-d:Z6�! {��B���
PB	\�ط'���s���]��b�e2��0�xf�� v�GV�%�EXTp_{�B��)��W�M�2��z��& ������d!��sy�3�E�':KQ���J�М�'���
ò֋�A�RT�;Cp�b��xF�a�Q�>/��=�䢘���((N�6r�=S��;*�������l ٓR$���7^�d����^�\y���^&Ir+9��)���<��b�3SJ	��ȪL����#|_��D��_	�:�@���Nn�Ў"������S�4�8t$�ՙ��^�Q����c����`��x���iv�i�����i�c";�8�ࠁ�Q,�
�GXKQ$ {z��w^��?�ɷ ��{�[y�8X��g>����bg����~b<6b��T��lt֠��M���q���(uf���{��k�Ӱ���e�P������u�gW�ah��`	����H(+���IT8�iz����_f(Vu�3�\�x>�n���y��8�雎��R���h��b�1ɏ_�&�j=2�o2�4&�mCwy3uq�@�����TuK;g4	@�Ō��pd�YN��e�n(S3��h�����V3�~E���yG�G���KbCG7'�5��+��N*�[�}�hY�U�R�*!�/˺
+Ʒ��󽑔cο������g_b�D�|O�+�p����"���}�O��[У�GRM�����O��Y��'&��#	j��G�˸)��(��g��h��l�	�w+I�}�e^v��&I_�g��%�O��`Jp���j���g��^I�2S�����U.��b�`:�L���P�#�#�Z�	��)��)Wս����T�W2Ԕ�lf�N���Z���#EO��e�,��-	��넚����)��[�BEo*�QH���Al�X_\�ѣ�,�Ŋ;V�T�P� ��Vo�V��3�h^m�Ԭ�|�5SL�Z�'Һ搜�&:|��E��_�7"h����*������}�
/H"L��i�~b�y)�^+�`;y�]%K�0+�	��z��7��3IJ��r�z��d��J��Py�G]�(DA�5\H�>h'c�Btư,:�Ya������hK�^oˢ��eb�	��dm���G��j�ӫ88���U�l��hGbɛmt��s��(aEJ�j��O�:�g�-1�(�k>���R���J>��խ��j=��O�	0�X�~69�Ȧ�<53��9��&%�M�db_�4�'�7�3�c�� i�?#B� _�k�#�:�����`i��T��;;�W�>#���h�4�^q���k�Dz��[	%yy*^t��$sͩ%Kg3i�"��:ޢ�D�r�r�"�B�T)����	@4E�~ʨ�M�ښE4m��ħ��ooǙ1��Դ��G��"ف�c�1������:Y��E�1K��?P��G����k�S�@OwEzգ��f�k�#j�>�nR��k�P��\��)j�4&���R]��A����`��\�	P�n����5��M�L��u�!��"�sQ4'�ͯ_4]F�}��k��·f�����_y�<Ҵߏɛl����F����Ƈ�"|������z�	� Ӌe�Ə���뱗鞵���ɣ&��h|]em��Kg�,�zt¨x3�sp�7QV���q���:O�	���Lm��g>bZ&)T����5J��)�L�.�a���E��(s,k�ȰB���R����N����E��72I��RY�qE�&
m4�� �"Au>E���˕)�#(-}��#nE>O������)W⋪����{bf�i[?�\[4��9&"��Uv�Xw��yr���D�.J8jŋ�X�?�η���t���鶶)���e�sC��+��#�&�,D�h��_~s�L�^�y˩0����z��L�t���"�tQ�#e�f���п2�9)���_��
�kY�(�>p�t�?�B�_.���=���D����M�?�E3�"d�����fՄ�J�����`AR���ch�?�7+Q~!?!+��@�o������7�����8�':�gz}k�,H�����k����Y�}�D��۱����>Z#{X�v^�
����.Qh�бDUtrO�����3W��^R�}uQ��9��d<�>�(,��&B�C����Jv��FV�?����E�M9z�?���PѓQ��i��#��;k�'E�J�.,C�����{����Ina�)� Uy��k����m@G��=a<:"�r� ꔔ����t���ef��;9���Y��Ʈ�(E��Q{�����D_�OH���\��}di��C��EY����m��Y�����>#�Li�Vu����]�≴�(TZ��.4��߹ag:�Z�%��\�����)�;�[յ��&�j�,�K��cZ|�~Ѥh"���
������'+� �l'K��3��)���A	���~D��"�Iղ���]}�>~'Zz�|���ě�	=���"X���w�
�O��q�68�L���o��5����H-������ `j�i93�w�����$�[�P��G��7�P� E����Ye2��U�w�􃆲^__�N�K(�|����i�/�x��Q����DT���YM�,�āW�R�!����2�|H<o!ԔO���������Rt-�����2c|���'=4�ږ'HP4�C��K�.�t���i����C�����,�T�z�j���;��uR��e�J�h�EƁ ���2Ņk�|=!�ϛ��g��x}D�Z�ohy��`�a�?-��U��4�Ð�ռ}ۼ�����l�����{V�Z�e5EsJFc��]4��Z��B�s%�
�}�#���s��0�TF�K:4����ͦn'�����I3����~b�sj�Oƶ��iY`��g��~O?6�[�����[7�U�l_�����ĮJq|Ôd�%%e��Y�s�O,6�?���٤9�<2�t�JZ�_{h��e��le#�pN��'l/��h+��)�C�Q���~q�4��D�8���t/|]��V.P�1�c�Z��xf���_��}��O�~'2Y��3�&]D��s�!�n� Q�ɒ�� �w�*�~�h���͘^֦-[��Tʿ/M@��R�f a�O�2⪫.Go"Z�ݟ!�
vL�!� o�K�n,ޑ��L~��9���:��0|~%ׄ{��Y̬�i/��V���,�m^�n�i�;H�ܡ��x+���`�+#9j'��	�^�%��R�֚dKaN�|ʊ�ɏ8��F��f�_�l�Ozդ������?I��f1�_?����4��z�IZ�E� �ct���ױ{�.s6���ڲ�@�3͞Ls����f�ɀ�SѶU�9Ȏ��b�މ�)Z-h���Aٰ��ѕ� q�׾~R{ I��;�p�A���X��~剕P<栁��22"�ƶC��M�̑^)��]q��f�A$�Nkg�9�O_� �%�ii�A�x�,��!����Q��I� َɶ����%k�m�N�t�B6��A�2���b���z�@�̴��

�fNw�L��Z�h9D+FHV��qR�W�9"��hӖ�̳��6֣���sJ~���_PGx�-B��#����5�|�^RAؿdV�ծ�Mz�@B��m�m�s��;3iVX�sJ���P�d�Y?5̼f��c���~�SE�JwO�aD;��s�����wj{�Ӭ��פ`N����;̃�[h���*�'nL��>b�Hr�T��a	��f���Z�Yǜ�gK~�ֆ-��ߌ�Ӝc{�-Qۨ+�a����0-Q��l,N�$)���U��	��q�7b.�v�V�zz	[$����u@PDѠD�����4o��0�b���Iԥ�F��N㱶�sc�_&�)�Ǝ ��N���?����.�	�t�����+I}�bQ���,��x�k]�Utޚ�8$ת�'M.�B���@)4���Qֱ�_j��)����5~w��s ߇T3H�RsU��5�W�����}ţU���\�`+�Gfj �Noǅ(i޼�~^�>f!]�X)��=ƴ���ƍ`$�y�`�9[��G��>-\[�����T��r����䊥�j��~U�QU�ʡ�B����1y�Y횷�&�b<�\v�	�<�i,�������uT��q�oޜWp�
ͥ�챿_>������4�̉�<-��*��U2�HEb&ddO�x
�i�w8��P���PRVk�h��9��hf#s���<����z>U���?��ivm�g�
�J ��<yfZG@����E{�+�RP�;b�};|&�:(5�1����q����n�n��㎙z\���ʓ�8
�ۉ��t��׋[1X�e`>��5չ�gɰm���	�tl�B*>�����go�#V<�������<�ʋ׈H(���~����b�W���`��W���Fl¼�\�=C�VK�m��,�Y0rUהV>?���m��BN��6{��/Z
�ͽ,�ydy�^����)��Л�5��8�a�?�K��p��Ճ�vl��h~?كsw��rPC���$��n+�ˀG�y˯�A�;�{�g45A���n�|�����s@$�bx�W��R��h	vPB�MtQ�r�{�zo�$�v���%o9]����A��nOU�Ie�� �������̻@,`�[�2�ɳG�ߞ���ۋ��yyv]l,�Ru͕�h��u$����ĎㄷT����~l�<�������VC㦦s�q0{ϓ]�Y=���Eu��T�����i�>�q>��TH&j.�ɥ~���yA$k.~]~�fֻ������]9�?e���(��5��(����]�\��:���ۅ�����_E/i�Ow.M�\*���6��O��:�;�L0�c����䏗��J[�����T=�4ц�ƾ�;��������P7^�MHx�T���1��.�l��v/
2����J��f���S��(S%g?��o�z�������H�n�s�)%��7S�K4T#�np���sCX\���煅l��|pÀ!�ր��k�杶U�q��s�@���CGD�A�|(
��O��ֵ�Z�����_���vxw1��E�q�9���
���4)�F@��Ed�eL
LkEA0,k=����KN�D�W�c���yS��|^��.`���B�L��8b�b�b�ے1E�c��ijϔ`�R�	c�qj��zŏz}�x���)���u�
FHحz��\a�^�!�V��r�[�u*V,���*�;�j�kt�ͺW--V�5���'��JQ��WT秼�+2�E o���v���ۭd+�q��AX�@������d����p:<+D��Z���q��j�R��l��W))Ca9���bP.Ƣ���|UsʚNmq�I�7�,J�V�4���//��-SK�z���[x�a��_�HH���k@���&�Q��-:ը�:*�� ?)�n�T�d��-�HL���L�
�%��{U�ա��W���DR�L1�x��$]Q�1��f�W��P��ٷ��TQk�&ܨh6,�Q�'����1��]Rm��:E�d�Q�_9M��o)(My�OH��%o�Uc(�A��sј�N�k4���hM���V��FZ�Sy!�Z(�sw�qY�����A� q�nJ���d����4ylm�d{3�I��g�A�	�&}@0��W�=�'�1����m��A��k�*|��(.B��VrW ��;��w񚋷������{.}@;�3�BKo�x��<3yNj���kwQ��C�?M�Lt�+��r5]�r����e��+�������9n˧��0R_i��j�η�>��ObH�{!7��p���mr�����G�D��]��E���u��ƌ���"�v�f��ܔa
�#P���6��~~�������z�W����Π~��Ք�Ib�r��;A=�
05�I4�p�ֽb�ːo�ĘX�ҎzJ���-���l��P�y��鷠�M��7����?�<ȔMBq{��T�eP���>b�\;��������ѽY�x����6'(�	�2�k��Br�������e�L��X$]?���AcG������������ȯ��s��{����]�4��H�V�K�~=�F��$yی�_�%�_$$ 1��_m�b�WI�ގ=L&iPt>b�1�*3�(Kߑ�+48o	z��dPֱ��w.��en�;�W�]:����F�a����g�,�hA3/}��������)r�P����R:j��3�������
�H��1h��q'h��+b*\J1�H��ko+f~\�H&�T&����	�^Ӊ�jm�>J�6����\�Gz�$9v��}�"/�
�3����������=�_%U��Z�,�� ���PWc/���aS��$�,T��{(�Or!�0u6!�F�'!�n�M�+�NR=�1�Cx�ҠU�R�|� (�V�i�w|�?�ݧA���M�	>����c�K�	�#�o��Ga;%�И}��x㋃�P��5Tu���8H�3���� �E�
E���r/�y����t�$IO��L�(�-:B�a��[qI�H�I��N@�<B�c*��V�
�,�2��C�N��@���9B��$��3��b������BE��i���D���\c����~�	�4��u��8���nm:��T�N���M��)�>0F1B����{�{�)X3q��Rք[ĮF4-��0����֣�"A_d�n�M]"ʰ�����B1h;7��Q{��tv�}PQ����R���9��%M#ҨWv��TR	[�W�	�@PA5�5��3e3w�\y��(�^!��[�r|��푶e��b��7d1(� E��ŰZ�]�r������m[����bL+F�wh�I&�d��w7q�2���G�_w4�Z�tP4�{�ɸ���f-�ă��=V���� �l������C�Q����KP��0��ɉ��P�nP�5�A)�V�x扆ʝ1Dh�I����zo�a��o:Õ���7�dd����J�C�-I hz�ѽ�L�0�� 	�, e��M�#�R�ߵ��� O�n����HL�3�|*(P�U��]t��IP7Q�]@�(]\P*���6����u�i����X����A[	�f:_dZ;^ۧAs�c��f�(P�vj�� �Ew��
�MmM�ff=B��QɅ(��~��Ak���e��L'p��든odؠA?Tڸ�5R��'x�G���A����4E��8��0�0��A輆>8�H0ꒊJ}�w^݂�T2��	�?b�{L������M+�p��RSjb��Ǆ��"��8L��*dl���o}O�V�FY��Jo���@ ��9�ul�f����8�y׷�H�ݎ�à|�h�`�K����L�e"�I��� �O��%��c��;�^�y�c��4�Xʾ�o��l��1�觩,,�"�(j�ϧ�q��߃��!��>�0���A���30;bkeJ�K�{�hӒ���?v�x[�w�xtf��ixƚV���,v�Ӎ��B�X��f���G%�~���ç8p%��pb�7��y�W���9=yN�>��N�v^ݝ�	��A�@�c���5�y}��W�JoеH��6C)�<�^�*6�PNh<'��R�'�:�	���DN������2�v�y��,���^u5&�d��+2�#f���_�v�������\�\m���,�8�/���s�&}�-�t|���A��k:���Ju�:i�)?��-��2Y�T� �CK ��g���lը��n?�G��Hy3�k�����4:�����}+]	(ko��b�ze��c�X��;E�;�T�ug�ul:@����t��F�JꏴWH�������֫dZ��~��X�ήn�]�f���6��[��%T]9Wwݠ�T@1ݱ�<��wP���㹺
A@���|�n�:�[�ʀj ����L��	&"s��-�t�l�&��JgN�%kB���.�%N1J�5=�N.<�P٘��o��.�~4kzyFr27�'Y��>|n	H��s8䥒�NcƤ�=�Ѫ���t��`�Ԫ�'B����wS"��6I�= �O�p�����y�<�q���ez��{�+��B�LM�_m���@%ED����^ī�K�>��s\�Q�9��-W-cp��f�a����pU۩���@�IT5^�|�{����;r�4�;f%`���B���3��ȃ������gO�3�V ��fַBI�𢝚9�(fIq|�� ��p��Vj�LD��)	��ռt|�ɶ$u��"�9��i\6J�c��}2�V#̤�+gR&ٝ�a�̪��0��%\q:�L����ѧ�\���_��7)+)���0��SC��P��fa� {z*����@%EE�:��	,cw���u��\���ZCY�/��8��fpTǩ�O�:ws_��pxe�j�8�C!4rk���� s6��~���J����T�_�T��jzZ\(0�{���0��3a�4�|�M�O��Zh*�^�z����}����A;�9C�� �����5�`(�K�'��d=���jo^�Qp�4�q��%do�$_�,wI��=_�&���#0����>��>���Gg{c����P��� ��?�|�p^���K��H�H)����{��$p����`�h��u�cuv� i�ų����Mda�F�������v"v��~n ���i�Y�D
� -rk��>" ���tޑ�\���2�;�B�fͼ&���Ҽ��DPUy�ڢp��5�����f�������>)�Zn<���#���5�Uz��|L�)�T�m����4���mz;P���%�h�;2�Q�� ��M�쒂$�&ԯ��OͲ�0��̎�p}������ K����#,Fߕ]����f,�Y�:f<a{�~y�pn�\d=J�����c�|p�s1�H ����g�M��n ,�L��aZ�S�L-�4��u���*��{�L9��zd@�e��1�Ș�X�C����7R*�G�<	�-\f*��ǫ�~��B+�Z>ڷ���c���f��\kj{����_-�[�T5���Ae@�T��5��,(c:����ZP��/��E"�7��/�����L|�X���*��]������G�W�p����-v� `�g�`�1�R�ioY}�M��^Ƈ���l�SȆ�н�w;�BW����S-�0󑾻j1�m���;R>S���?��b���]s���O�n�8�S:�J�X��
�,��ס.��u�И-Em�ӟ�?��ܰ�em����xA�5!5K@^Qx;���`��m�p����Q�W �Rl�*�؏�{w���ex��eh��#U�B�qm���	*n<�
�;	�Y��]I����Y�+��=E&���i��4�u�~V�H>��~�s���[���m��3�L�&i��(���nHPdpb��Ϛ,J3~��O��iH�J�v������n&����}5?�>I��?��Y�Wta��0O+C�;]��CkS�	܀-^nsI7�xwle�gJ������2�t)M��t��i�ko9������79eC	#�<	SS,�=ӭ�j�:l�;�J��\�H�>������:�=�,$Kc	�MMgZ��֟����Tk��P��S��`,��	d��a���(�A�";.�K��������6�M��os{Qҋޕ�������#�D�m>Z�Tj�D_x��R���ff��g��$6�6z2���JT�K���.1���>o�#��cw�8|J[���p3+����$��{̨Ix��$Oi����˥b��c"��\��AJ*e]��^�<h&�J�{L����[��+�q^%��y� ��s��>K�=���G߳ �� ��)Х�Y�ĵn遀�F�UEh	=�<[��*��P���Z�x�V6�(8J�ݨ�T@r�~p)l�w5�j���2�;S�fr��r���%'���8f�y����2�K4U���7�8X��:�
��=���4+�4]\���N�Dвq쭠>�q���7�����������"���od��tu����]b�/�������x�w[v���B<f}�<�	)�bNҊu�ќ�#?��O.�ɳ%4l��5h��AL�y��T��ξ'�I��+�&����b��J�뭒�ؠ+�O���������r���.��+�\��	�p�U�v�Q�&oe� J��x��ͥ�ԍ!���`)dGF�+	�c5L`�����P��]�>3��I�m�9�)*kL9�/�le��Х;d��O!T���Cʚ��*ye��.����؏��Ӏ�p%�{�?\iG��h�7�d��]՛���:���E��--:�W� у,�ą�Bǻ\3LRY�z�e�T��%�4�F��d:�	/M_��"G���S�"z��,��oz�Q����b��B���v����k[��1jr�nU��#C%P�i���v�l8���3�h��O��}�Z-hP�f�zeF}@6[Z�x��5�OeA�?�
���x �M( s&���I�uYJw���=wd��0i�sC)i���v/N�1DA�T�t, V�Hٳ����!E��aV��&:O@���MEߢ�RN���Yǵ�>���i؊��k���e.�ڷ�ٱ��巔RiR��:����јUK�ӹ�#��v`�V���'��un�pY}���l{Ŭ��7�M����1�v�/6!y�.هyK��j�)��,{b�^��k)��)��E\�
��0Pcy����<{ �w�,Ͱ~_�����iVu���|\�Y�I?�lS�.ţ��wXi�;5$��eS#q[��nG���(��όap��D���5�+I}���܈~����sXQ&�����U�ۀ�H�k��R_��M�V�@K#^V�٢�ܖ�49�Ĺ&XTd�؜kl��m�EB郖N��U�� ��sY�a���C�m����d�YڋG����[���%�649E쓱ۑ�(�`�]X�̓�ST�'�k��!��N����i/V�n�Ƕ)V���굤̠�OTQ"Õ�X��pZ���kY|p<(<��ҏR�
�/,�/����̩�5�y���x�OM�7�:�5�w�*���;�S�1�:8��O�Z