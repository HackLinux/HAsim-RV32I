��o]�����7e��u��Y�'��{����U��r��b�Y���n����!ae�1f�����c�^�;�\���Z�b_��0�
J�����V���,�#�ȩa��*~"����<x��~�/xT�2�?��M�܇�[��=�^�_|�Q÷���2P)HѨ<�[�h�5<qAz��1֙�>�}���Wj+7��D'Eh���s>�&��ow�p���B�2c}º{3���;�l�į���C��$�V^�-m�=�Evo�/g�����r�v�#�|5��g��+I��S��?�*	����ca�G��P8/����6~�Qx���=� �M�k�3_��@ IX�g{��R�4�ƈnޖ 猢�h㿬R.��*i�����������ސą��ƭ�M~��J��Z��\iF�E�0NK�(�.�0{�
�=,����``$�;�	

h^{7#oG���	{�h0b�Yv���m�P�F����$#Q�t4\LîQ���5��1��@� 2�i<P�q,=�\������^�<�gSy%!��{��W\�ho%�K'
g�yAkO2�l*[�_��B�U�V)@�����]E�{�hgU#�c�h��ޏ�ޢwU����Z���*�'�3xZ&tJ�@,����WLl:-(ɛZ�!�$�=$��v�6���t8b`�M�iO�o\w PI�Ӈk?��M8J�~�)���{��r=3x���&E�U$b)dP0h���ȣ����p��cL�GVZn(J��^&i�HIV  ��\Y��\�-�굧��ߕ��%a-)-���,75�%H^� �T ��Jܗr�t��)��WO� ]K'ҟ+4��-��'(��B���b_��i��pv�����Uupj��MDw��U}ژ�_M�VW�9IR�9 |d�vV��d�_��E���FY9�&(�X�t����m�|seHre���v���`�����]F?_���3��*�� :,2���e���
5�!��%$3GS1�`o|�C�"����m��}a*$l����Ǝ�D�9�*xD���C���{���a!Q��	z�v��w����4� �T���te1f6N�����sEf[�A.��᤭!�{E�ޏ�i*�����i���x�Aa���o9�r�7V̷������w�쁎:0�%��$tdI���(��i�C�N%�
� �=��D��P�����|��X�6�2cW����D���m�"1$�����y	���Z6���:�݊���nS<0M�%�́�����>�e���}�Q�DV�3���i@Bf�$-E鄛b+H�C��Di�-��������O,�,�u�t�uSO۝b�H{c�X�������?�����m1Cb�Q���7��"���'8�8K��Ο��Q�T�C�s��������f������m|J�&x6sGY�;I�'�#6�=�����U¹� 7�Z��Y��zv����2��fu���u)3}�?6�_��L��:6��(�xP����P�e*���T�~{t,j����_R)�S]��@�3�p�TP��y�	)�6h����I��f��(���v)U���/�1�7�n�3���$K�\�{�g�E�NK�q����U�>Xc��ժG��9w�ۚ�|�a�'q3ݚ:����a�ɹ�G;Ձ�_
|��������@�5��?b�ĭ�d��ې���h�M������8*���L�t�%u���	0: �^B��S�In��	�NL��h�[����#u��G�M�u�1-�,O����1�UůxN#�q�iǍ�Z�$,=x��9���9�zmJqT?��튋���l?����%-
F3��\�H��-jKP�b}E&ȹT/�n��X�����9��r�кE����&ŝ��])�`�6�t��+��Q'^V��ڲM$�߽ywUg{�sA�Es<�,F���F�`����#�{��/��D ���E6����?�QL���%C�=t7�;m�*�TXdl<��g�n���NpbM.vC99E�����S,���J#Ƹ��f0 @En�����]S��8�r��|�6���#���i^G�|h�x��X�	�z��5��Y�c�q���{B7�o&8q�F��K@ ��]��$?�ُ�TV{�U�h�cE)!��T�:M."œ��?�!	C�<G3�)5�>��!+X����'�K�M�,�����/�Q��r|�)8#-t/���A_�{�I�����	�\*%O��-I��aށ�Z���s�3\FґE�Q�l�L`�@���KRSK"T��zj���j�h�i�U[� ?�����~� �wo�:c�rUȯ��M�	�❉����:�����|03�����	$�f����ד#��DӱB�㶥s'�������� �
f���`�*�Hhh|)������r`�B��}�y����^J��ʰ/��O���S%N���h&*t�M���T�ߔ��
a8���vB��Tɧ�kQul�(k�į�2n�L?���2F���YX\['�#�Q������;�ŮX���^�"Ȃ�2��uv?�����&�Xf�=4�x���� �d�!��u�2�v�.�V���O"�eo�շ��2�����V�3��B7���l���H|�M�^Vxɝ�{Wl������9º�8V1����L	�