g�r��_r��F'9n�Fڋ=���Q;Xl�)�h=�u�@Ol�����z���B<�pGzI�G]��{���\͞�:�{4v�-��g̕�����r��z�������A� �?�k�N������;���l��"ڞu�X;u׷!<�$-�y��h�:)��VƔ�OA�EB�����D��@��?�7�L[`�H-�Ei�dJv���x#?D�D_Izc���Sp'�+ж<@����:���I;j&��;M=�&��#���x��w�b���M�&� ��<�o�g��2��؟�-�ӛ����#|D�2Q��~�3�g�������[�7)�I`��⒅�|���c7'�C��,�7!B|���ƞ�����Sc����e{d�K�@�kP�x�G={�Je���~�?9"���i�.@��0'��I����L]=.���{��g��b1�H���ޯ������j��F��⬂��p� ���O�n�Zҍ+�6
��e�/\d��H��BK�I��C��K�G�l�� �FL=�J���>�4J��jwX��B�Ԧ.�t�}���P	��M�x���'|�c��h��!�A������p�v�,��MyaISj2���ha~?[1>�HH��~�/�1��nHx�j�Ҹ�hUT���LϬ�< z/��+� Ȣ{�.:qc��}DP\�ċ�ջ�Hj����w;L��7IK�c<��������p���7@fggjG%�1PO%��E�tZ�a6Wb��SE�GdyFʣS�_	�-���q�LK���'�����������ȏ��ι$�#[�6�O��Ō���$�AD��uOWݨk���B�ʔy��}��D��'k<g?���L�2�!G�k�����x_+6A�0�j�������c��c�&gU�΋�%SU��+4��,Z��c��w��K���cX�D*�r޹��Xܠ�{��bg��a�7��#�����c�zO���i�om�ڌ��N��ӫ�E\�*3�P7&&k[�LCs-u,�⫷K3~���90���(W:�ec�Ϛ�6�6�P�	��j����Z��T����3��⌖���\��("�m��H�윀ն���_��@&�#��H��x������j���lر�"�&��L2��ݛ�
��f��zl��"��,"�����B'2IW��/�v�"� q�[o�����:^f�"�����O����t*��"�A�Y�&2�QL�)������7M� ��}�bp������.(P�!HsA���>�)�󒠊��諲��~����ݠ|���mBJ��#5����4��k�ݢ��`���T�����'x<�����Q8~�fn�Ґc��k�Z�"�p�$�"z��$��&HZ6�&��Aw��Z�WB�_�R&���w�A�!]��z��X��6s�H���U����rA4e7�*p&�]�kB(lF_Wڿexj�͑��V�̎�S��-d����.G��H�ź@�ݔ��9��)�&j�K'�S����ơo��%ݷ�F�Ԥv1
��rḇ Ӈ����Ld�r7�	lr+b����N[�ͪ��-��8u��D{Un�ٞ���rz��>Ҽ���zh�5ޤS�O�U9�`����ySR��������&xF�L���8�x0[���v�e�	�:|0���&y��zq�%k��>�|��2rS�r\)7u��	��w��a-��h �w�>L��r�V0Yw?���XC�	+a����1������0�D���d�2���e���� �5�$��:�0�r���Qm��yR�c��am�kmw~=0N;`+�z����jC b����� �q0��Բ�/�Wы0Hxvѭd��P�*�G� ;�p��^Z	�<�2�0p����q�%��,b�0�	���}���+�����5��rm嫚�vK*�;�'=h����$QYdXvᗤ�U�I�-���脯8 D+�+'��ɇ����$L��X��j��=��E�`*�B��|���^W;���T������6ͪ�뛔�B4Q�K[B�͡q��Hk�����B�����h��'���7��1
�R���,��A&:$�m���U�ޒ��]�fc��� �LkeO��������:D��3r
�T|fi��]c�e޵�2�u���ތˆ����Nxe4!��s�8|���Z���IE���P��?����{I"�a�ڎ��<�.�X�`\�	�=QgB΄�IHY��b�xY��o��w����X�y���^F�߆��T����yF�>�KO�Q�0�4��Nhw���f�$�!��-�g{� ��>Fl��TNF����`�ݻY^�Wh�[����K���i���AXE�4��S�fH�53�>|�#�m�Y�[*{Q[�'6�_�7�^c�t������I�ɼ��(BM��8�LnVo^��^!6��5I��|w{L�S�X���Sj$��-��݊���� N� ���S�0�R�;�R��|�ͽ3~�ѷ�A�4Qi� � �5.�[��'B&Q~�d��!��p�+�W��Ȅ�Q}�u�V�b���d�}:��D�2�&���Á�1gh�c`5���h�4{~hF>+�'GG�	��F�������9�?d�bh�\S��^���َ]/t��+�O0Hw�\�Z'i��_=&jU�*���Ƹ�ʮQ�v����d��3�o�0�8&��ޜb���/>c��/��̶�"��х�^�J1-�}�i�KK%-5U�@!���j���O��m8�����pn�o ,z7/	o��6�8$�m�$�#˶�J0�]o��s��쫲e	ʠ�=�|����F�l�����Ym�c�k���P�ҚPd���G314D����T���0	ˊ��$�f	{�	��l���k{[I�}��0���JL��ZFi2�Jw��|�w���׎!m�J�3U�P�2�3-X"���%t��I�n�r����?�%4;jh|�6�s�E���"�gKk�	��(v�j�w�������,����X�O�c$��4��Tc�75s�*j��
6������]��� ��uy:�n?j�w# ��?���s3_���9��@�j���V\oly�,]]����obeo3?���y�Pn��@Z��@��v,����o�:5@�j������QϪ��o(/��It�~S�L�a@c�_��Xr&Q}i}�!��7C?�b��O�@e�Y;�� \���)���ԭn��.�[����n. ����1�l�N�TJ|v�����ZɊ�HN��2���-���ռV�J�_�V����8���y�k@]Ę2�YXx/?���r.�oU������Q"�!F���+���?��S x��ޒ�W5���+&�e��uJkR&@���26�?9Ir��j�럪 l+s3�L7Έ)g������Z�����j�3�i[/�3��ڇ���f��@�[�j�"��o�$Gb�3��Ё�j���uB��>B��LX��_�*�us�ON(T�?#�i�� ~����mZm|/`��������Z|(F��������8�j���S��X����]�کJ�]�J�BȡsMV"e�df�����[3v�W��<<�=o/�n��<�'#Z�u��V�2��_��)�?�T����5YW��I>�b�5j�����_���U���U��m�L��I	>�]I��7#j?�xW(�hy��01�6��	槌J����fH�J p�*��Υ�7���g�u2a��L�Me��@�
�̑vA6%<N9|�������{^���9���os�r��(Q�Z^`ԍm���IUD?��S�"o���?)�Q���J^j�B	��b��y�*���ݝ���1='�x�!�I�_P1�X�8��>��?Y��K�Pg~PaU���]h5��;?��6x)�����Ubc!y}��fc}�`im�u������Imfl��S���ș8���
���?J���sH�(�հg�Wg��]�>�̡�B��^���x�%�聾���%?ul�M6v��=�e��
��u�%�ԠTQ�W,����N1��iӅ^�99=����Q����WR�w�p?�c�h�č��f��v�3��� ��ß̬�ù<�9��s�Y�2��M.L�B��2�Pq�Aqes�c'��,�Yӕ��w�?7����Ru�./�^y�E9�`���P#����*Z-r:���u��|�I����K�-pR�1`6��}����ʁ�a�Զ��/��5�E7١DZ��ە�x��W%�Bk�n�&���`�0�:�,C!-�yl_i�遝+���i�LOL�p��0�чEul���.�h�<��M.���e��Y��H�C���N�p�齢����^�"�Dӏ�뗖��6�����ச���φ��Z��X�!w��f!Q�����"��-��6�@�<u�!(���|#�=:��#����|��