��������������ή���ݾ�����������ΰ��������������������������������������������������������������������������������ν������������������������������������������������������������������������������������������������������������������������������ӳ�����������ӹ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӻ������ӷ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""&P2K3PR3K3RKRK32200202000200.0-00E00-0----,$,#!#!""!#.KPKWX\\ee|������������������������������������ͱ�ͯ���������������|||qe^^^[WWWRRWR3R5WWWWWW\\\x|^|�����������������������������������������ͱ����������������������������������������������������������н��ܽ�����ݱ���������θ̯��������������������������������������������������������������������������������������������������������������������������������������ӹ������ӹ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӻ�������ӻ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""""P2PR2R2R3RKR3K22302220.2P220.00.000E0,.----#!###"",$.KPSWWX\ee|}������������̱�ΰ����������������ν��α��������������~�||~^^e^\WTWWWWWRWRWTWWWXW\\^^e^||~�����������������ܽ����������������ܽ��ΰ����������������������������������������������������ѽ�н���������������������α����������������������������������������������������������������������������������������������������������������������������������������ӹӹ���ӷ��Ӷ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӻ������ӻӹ�ӹ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""RP2R2R222R3KR32P2R2R0.22PR2.0020.00-----,---####!"#""##&.PKRQWUX^^e���������������������������������ݱ��ܱͯ�������������~|^^|^ee^\WWW\RWW3WWUYWWW\\\\v^x^^|�����������������������������������������ܱ�����������������������������������������������������α��ܽݽ��������������α��������������������������������������������������������������������������������������������������������������������������������������ӷ��ӹ�ӻ��ӹ�Ӷ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӹ�����������Ӿӷ����ӷ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""PP5.2R223PK3PR5K3P5222P322R2K0000.-0,-,---#-#,!!#!#"",--.IPK3SWX\^e|�������������������������������������Ͱ�������������~x|^x^^^^\^\WUWUW3WTWWW\\\[\\\\\^^x||���������������������������������������ܽ��μ����������������������������������������������������������������������α̰������������������������������������������������������������������������������������������������������������������������������������ӹ���ӹ����ӹӹ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӾӶ��ӹ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""TP0P22R2RK3K3PR2R23020P2P222KK020-,-0-0$-,$,##!###"""#-P.2KPWW\Zeee���������������α������������������ѱ���������������|x|x|xe^Z\\U\[WWWRWRWTWSWYv\^\\[^x|�����������������������������������������ܱΰμ��������������������������������������������������������������������бή�б�����������������������������������������������������������������������������������������������������������������������������������������ӹ�ӹӹӹ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӿ������ӹ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������!"""""""!T002R001R3K2K2222R020022202.0020-0-,-#---,$,####"""""#-2-0K3KRR\e^eq�|~����������������̰��ί����ѽή�α��������������|�x^\\xq\\Z\RWWWW3R2RWRWWU\W^\[\^\v\x���������������������������������������ܰ��μ����������������������������������������������������нα������������ΰ�����̯�����������������������������������������������������������������������������������������������������������������������������������������ӹ���ӹ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������黹���ѷ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""""""5P022P202R22K2022R22R21.222.0002-,0--,-,-###"!#!#""$#-.0.PKWKW[\e^e|x|���������������Ѱ�������ܶα������������������~^�x|Z^^\^U\WWWWWW[W3RTRWU\WW\\\\\^^x||����������������������������������ݽ�����ܱͼ���������������������������������������������������������ܱ������������̱����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӹ�ӹ��ӻ��ӹ�Ӿ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""""P00P223P22R222.022R2222202022.-0&0,--,0-,$#,!",!!"##-0-2PRWS\\^eeqe|����������������˰�������αѮ���������������|�|x~^^xx^\\\\WKRWWWTWW3RWRWW\WW\[\^v^|�|����������������ν�ݱ����������������������ͼ�����������������������������������������������������������α�νѱ��ͮ���̮������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӻӻ�����Ӿӹ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""""1P0102P3P223R.0222P22.0001.000,-/-,-0--,-,$#!!"!"###.00.KWWUX\^|e^e~����������������ˮ����̱�α���������������~||~qx^^^^\\\\\WRR3WWPRR3PRRWTRWR[\]\\x|~|�������������������ܱ��������������������Ͱ��������������������������������������������������������ͯ���Ͱ��ͱ��˨����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӹ���ӹ����Ӹ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""""P2002222.0R22P2.013000./221.0,,0-/---,-#-,####!"!"""#!$,-0K2KWRXZ^^e|q|������������������������������������������|^x�xx^^Y\U\YU[ZRR2RWR252RTWTWRW3T\]\^x^|q�������������������ܰ����������������ͽ��ͮ���������������������������������������������������������ͮ������ͮ�����������������������~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ӹ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""&P1022022.22.3P&0.000/.0,0,,,&,-0,,-,-#-###-"!""#,---0K2SRWWZ\ex^^||�������������������������������������~|x|x^|\x^\\\[WWWWWW3PK3R22R23P3PRRRWW[\^^^||�����������������Ͱ������������������ͱ��˖������������������������������������������������������������������������������������������|�||^^\\WRWWWWXWWSWWWXXUWKRSRS3KRR2K2K30KKKKRKKLKGKKIJIEEEIIEEIGIEIGIIJLLHLMLLLMLVMVOLJMLVMLSMLMSLS`Vf�}�������������������������������������������}dccXURWQWTWRWRWWW\ZW\XZXU\Z\URWRWWRRW3PR2R2P3R.R3K2RK3K2RK22.02220222220P22R3RRWRWWWRWWZXWRWRWWWW[W3UW7WP\WTW[WWRWWSRWWK3.PR220220201002222P30RK3K3KW2R.2R3RP3RR3TK5WRW\W[YWW\W\WW\\WRRRWWR2WR3PR230R23PR3P322R2K2K00.2P20022022222R3WUSWSWXWXW\XWWSWZXWUUWW\U^}|�������������ӷ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""""P5R22222220K3Q220222202220000000000,--,,$,###"##""#,0.P.0RRWWXZ^||ex|����������������������������������������x�x�|~|\^Y\\WWW\UWRR3KRR3RWR3R3RW[\\x\\xe|�|������������������������������������ܽ�ܱα����������������������������������������������������������������������������������������������xx\^\v\^UX]X\XWZX\^XURWWWWWSWSRRKRKWQWS2KKKKKKLKLLK.IILIIKJJKIIJJLSMSLLMLMML_M`V_VLV_VOV`V_V_Odd������������������������������������������������|fvccU\XWWW\U^\^^U\Z\\\ZZ^^X\WUR\WWWWWWR5W3RWWRR2RK3K3RKWR22R23PK3R2RR52RWW[WWWWUWWWZ\Z\\UW\U\U[\v\W\W[W\\\\WWWWWWWWXWWR3K3RR2R3P3022R2R3R2K3R23KWWSWR3PWWTWWWUWTWWWT\\^]U\\\YU\Z^c\[RWWUWWWWWWR5R3TWWR2R3KR2K3RWK3P2K323R2RR23PRWWWX\RZXXZXZX^c\\W\W\\\\c^e^|���������ӹ��ӻ�Ӹ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""""1P2R2000.0.2K3K30000220220,,0,-0.0,-,#$#,$,##!##""!,0I00.2KRRZc^e|�q||�������������������������������������|x|^x^|x\UWWRWWWWWWWR3R2R3RRTR3P3RRW\^v\\^^^e��������������ΰ���������������������ͱ��μ���������������������������������������������������������������������������������������������~^^\]\\^UWWWWWSZXZX\\SRWSWXWRWW2K3KRSRSK2KI.IKLKLLKGIIGILLILKIIIGJLSLMLLLJMJ`M_`VOVLM_V_V_`VX_df������������������������������������������������}fcec\cUUWWWW\\v^U\WWWW\c\e\YUWWS[X\TWWR2R2WRWW3K22PKK3KWKR2222R2RR3R30R2RRTWWRW3PWWX\\\\\[WW\\^]\\\7WWWU\\[WWWR3RSWSWWWKR22R3RR2R00122RR3P2K222.WW3WW3RR3UWWW\WT3TWW\\\\[WWWUW\\\^U^WWWW[\WWUR3P3PRRWW5222022KRKR3P222R2RRW3R23PRWS\WWRWRSWXZc^X^U\\[\^^e||e|�����ѷ��������ӹӸ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""""PP23220.0,02.R0220200020201-,0-00.0-#,####,#!#"#""##-.0E002K2RWZZ^^|exe|������������������������������������xxx^|xx|\\RWRR3WSRRW3K22R3R2R3R2RWW[\^^^\\x^e|�������������α���������ܽ���������ܱͮ�Ͱ�������������������������������������������������������������������������������������������~���x|^^x^|^UWUWURXZXZX^SWRSWWWSWWKRKKXSRXLKKKIIKJKLIKLIEIIJKKLJJKJLLLVOSLLLLMJV_V`V`VLVV_OV`___df��������������������������������������������������|}|c\^cUTW\\^^^e\\W\UWX^Z^\^ZWWWW\WUWWR5RRWTWWW32K202KRK3RR222KR32RR5P3RRWW\WWWRWTRZ\W\\^WUW[\\Y\\]W[WW^\^\\WRWRRWWWWWWW3K2RR3P3R2222R3RWRK222P2WRWWWWWR3RUW[\W\TWWW^\^^\WWUWW\\\ZU^UWUW[UWWWWR5R3RUWWW3P2202KR3KR3P20KR3RRR3PR3RWW\XWWSRWR\X\\Z\\WW\\^X||�}����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""""PR3R220200.02.02220022202000,.0K00.-,##",#!"#!"""##&.00.022RKWWZ\Zx^|^������������������������������������|x|x^�x|x\\WWT3PR3RK3R2R2KR3P3RR3RWW^\^^^\^x^||�����������˰�ͱ�ν����������ܽݽ�ݽа��Ͱ������������������������������������������������������������������������������������������������||~�||^^\\\UXWZX\UZ\XWWX\WXWSRWS3XXXSXRKKKKIKLKILKKIIKSHKLKLIHLS_V_VOLSMSMNVVOV`V_V_`cV`cbcf����������������������������������������������������}}|c^\vX\\^exee^\\\\\\X\\U\^\WWZ\[WWWWWRW\WWWXR2R3P2K3KK3RP3P3RRRR3R3RR[ZUY\\RW[WUWZ\\[^Y\\\\v\^\Y\]\\x^^x^WWUTWRWWWR3WR3RRR3RR3P2R3RWWWRR23R2R2RR3RWWWWT\WW\[\[YU\x^|^^\\\\[Z\Z\U^\[W\W\[WWUWRT3\WW\RR22R2K2RK2R3R22RR3RW3WRRWW\\\X\WWUUWXZ\\X^v\^\^|^}�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""RP2P22000.00.0002220.R220.,0./.00.&-,#-#!"#!##!"""--,.0--2K2R3WSW\^^|^������~�����������������������������|xx^^xx^^\URRW2R3RK2RKR3P3WRWR52RWRW\\\^^\\x|^|�����������̰�����������ݰ�ܽ���ѱ���α��ͼ�����������������������������������������������������������������������������������������������|�|��||x\\\\\XZ\\R^U^X\\\Z\WWSWRSZXSWSKKKKKKKIKIKHSKHLSLSLLKLLLM_SOVVLMXMMLaVVM_`c``dfdffdf��������������������������������������������������������}|ecv\\^xe^|\\\^\U\^\\U^\^\\\^\\\WWWWW[\WWW3R3PR2K3R2K3RRR3WWRW3RRWRW[\\\WWW[WWW^W\W^\^\^^x^x\\\^Y\xx\^\\WWWWWWWWRWWWR3WUWR3R2R3PWRW3WR22R3K3WR3RW\WW\]\\\\W\[\\|^^^^\\]U\U\\\W\\\\\v^\YWWRWRWUWWWWR2RR32KR22R2RR3RWWTWR3RWR\U\\\[WWUW\WZU\\^^ee|�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""PP22000.0-/202.222P022222.000.000,-,#!####"##!#!#"""!#,$,-.,-2.PKWXW\^^^^||�����������������������~����~����~^||x^xx\\WRR3R2P2RK3P3K322WRK3R3WUWWY[\\U\W^^^||�����������̰����������ͱ������ܱ���ή�α��������������������������������������������������������������������������������������������������|��||q\^^\U\Z\^X^^X\\\^\X\XXYXWXWSSRKKKKKKILLKLLLLKLSLMSLL_SLV_LVOSNLVLMVV`V_d```cffflf������������������������������������������������������������}^||e^ex^cx\\\\\vX^cUx^Zc\v^^\\W\\\W\\WWRR2K3P2KR3PWRR3RRWWWTRWWYWU\WWYUW3UWW\\\^Xx^^^v^|x^^^xx^\|x\\\[WWWRWWUWW\WWWRWUWWWKRWW2WWRR3R22R2R2WWWRZWUW\\]\^\]\x^Zxx^^v\W\\U\v^^U|\^\\\x\v\W\\\W[WWRRR22R22R3K3RRRR2RWWWTWWW\WW]UWXWWW[WWU\^c\|||}|�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""""""""""RP02001-02.K2R02R2.2.P0002.R.020-,-,,#"#,##!##!!,##""""!#,--#-..0RRWUX\\^^ex�x�~����������������������������|�||�||\x\\[WR2RRPW3RRR3RR22R3P3PWRW[WU\W\\[X]\^|��������������ͱ����������������������α�ͮ�������������������������������������������������������������������������������������������������������|^^^^exe|^^^e^^c^^\\Z\^c\X\XRWSK3JKSKSSSLSSLLLLSLLSOV____VV_SMSML_```d`cdbddfffl}����������������������������������������������������������������||||^^evc\^^^e|~|vex^^^^^\\^\^^\\^WUWWR3PR3RWWRWRWWWRWUWRW\Y\\\\]\\W[W\T\^^^|x^x|^^^xxx|xe�|x^�x^^[\\TW\\^\\[\\WWWW[WRWWW\WW\RRWR5R3RKWW\U\W[\\\YvZ^]^^|^|^|xx^\v\\\^|^|ev^xx^Y^x\\v\\^\\\[WURR5RPRRWWWWRWWRWWWTWR\[\ZU\\W\[UWWU\\x^x|^|��������������ӯ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������""PK0000.0,.202P.P23P22P220000.00.&-,#-#####!!#!!!""""##-#-,--02KRRWW\^^^|^�||~��������~���|�������������~�x|ex^x\^^WWRRW22RR2RR2R3KR3PR3PR2RWRWW\W[W\\\\v||��������������������ܱ����˰�������ν�ͱͰ�������������������������������������������������������������������������������������������������������~||^x||^|^||^||xe^^^\c\^\X^UXSRRLK3SLSRLSLSS_LXSOSL_L__V_cVVVSVVL_```dddffl��}���������������������������������������������������������������������~�|ev^^^^\^|xcx^||||x|^^^^^\^^U^\WWTRWRRRWWRWWWWWUWW[\WW\W\[\\^\U[\\[W\x^^xe^||��|x�xx|x|�|x||^\\\\[\]\\\\\\\\\\[\[WWUWW[WWUWR2RRR5WWWU[ZU\^^x^^x^xq^x|x||x^^v^^\v|^x|x^|ex|xxx^^\\^v\v\\WRRWTK3RWRWRWWWW\WWWWWW\T\\\]\\U\U]UU\^^|^||����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������!""""P2200000.00.0P.0K02202220P0.000.--,-,$##"#!#!"#"""""###-,--,.0PKRRWW\^\\xx�x���|�������|��~�|���|����||��~x^x^\\v\UWRRR2P3P22K2R2K522R2R3RRRWRW\XWU\[\\^xe||���������������ͱ�ѱ�ͱ�ΰ�̱�αα�ή�����������������������������������������������������������������������������������������������������������||�||e|e|e|q||e^xe^^^e\c\^_\SWSWLRLRLSLSLSS_LSS_SV_V_V__``____V__`_ddddff�lf�������������������������������������������������������������������������|||^|^x|^^||e|e||x^|x^^^^^\^\\\UWWWWRTWRWSWWW\[WWUYU[\\\\\v^c\\\\\\\^\^x|e||~|~|�~��~|~|~�|^x^^^\U^\U\\\\\\vWW\\[\WUWWW\WWWWRWRRWRWW\\[Z\x\^^xx^|x|x|q�||xx|x^^^^e^|x|e�xxx|xx^^^\^\\\\WWWRWRWRWRWWRWW\TWW\\[\\\U\\^\^\\U\^ve^e|�|����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""""P20K02.000.00.00.2P200222020.00.0,--,,##!#!!!!""""###-#--0-0.0ER3KWW^\\\x|||~|~�|��|��~�|�||||�|�|~�qxx�|xx^v\\\\UWWR3R2K2K0K0222R222PWRPWRRWUW\\\\\\^^^c||����������ˮ���������α�б̯�������ͮ���������������������������������������������������������������������������������������������������������������||||�|||�|^^||qee^^^\c\XcZXSWSSSKLSLSNS_SLXV_______`dc`d`cc``c``hfffl������������������������������������������������������������������������������|��||eee||e|x|�xex||x|x^^\|^\\\[\UWWSRWWRWWW\WW[\\\\v\\^\|^^^^^v|^^^^exx�x��|~�����~��|��|~^x^x^\\\X^\\\\^\[\\Y\[\U\W\[U\WWUWTWWWUYU\\^^xv^x�||~|~||�|��||~|||^ex|^�x|�xxq||xxx^^\^^UvYUWUWWRWRWRWWW\WRW\]\\\v\\^^^^^^^xe^ee|}������������������ѷѶ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""RP.220K2P.0E00.00.2200.P.0020-02---,--,$###!#"""""##,$,-.0.&.P223WW\\\\\x^|||x���||�|���||||||^�||�x^^^|^^^\\\^UWWRWRWK3020K00223P20.R2R3RRR\\U\\\^^e^^c||���������������̱�αα��б�����������������������������������������������������������������|��������������������������������������������������������|�|��|�|��~e^|}xee^e^ec\X\XcXXSSLSLSSSS_XSL___V__`_ddc`cdfdfd``fdff�������������������������������������������������������������������������������������|||||||||�||^|~|^^^^x|v\Z\\^\XUWSWWWRW\\UWW[^\\\^\^xev^x^||^|^^eq|x|~���|~�����|�~��|~||||e^\\^\\\\^^^UW[\\\\U\\\\U\W\\[\\WW\\\[Z^xq^\x|�~|�|����|�|���~|e|||^�||�~^^||xxx^^^x^\\\\]\\URSWWRWWW\\[WW\^\\\\^^|^^^e||||}|�������������������ѷ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""""P202-2KP.00-00.P.0200,.00000-0.0-,-,-,-!#!!!""""####$&.--0-2PKW3YWW[\\^^x|e||~�|x|||�||^e|^^�xqx^\\\^^v\\U\]UWRR3RWKK2-2I022.2000.2KR2R3UW\WWWU\^exe^e||����������������б������α�����������������������������������������������������������������|����~���������������������������������������������������|��|��|��|^^e|}||c^e|cc\S\cXXXSSLSSXSS_LVSS___d__dcddd`ddlkfdddlfl��������������������������������������������������������������������������������������|}|||�r��xx^e||||^|^|^^\UZ\^\\URSWW\\W[WWW\U]^^^^x||ve^^||�|ex^|||����~||�����|���|�|^|�||x^\^\v^\^]\[W\\\]U\\\\\[WW\\\\\UW\\\^^^x^x\^||��|������||����~|||||��|~^x^x|q|^exx�^\\W\\^\WWWWWWWYUYWWTW\\^\^\x|xx|cx|���}|�������������������ѷ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"P02P2E20K20.0-0.202.000.200000.0--,-,,-!"!#""""####---.-,.E0RRRWWWWY\^^^x^x|�^|�|x|��eq^c^|x^|^Y^\]^^\\U\UWWRWRK2RK300.0-2202.022K2RKRRRW[S\\W\\exZ^e^|����������������ή�����α������������������������������������������������������������������|�����������������������������������������������������������������|�|���|||e||c^c^__cXcLSSLXXVX_LX_X_dc_dcdfdcffbfk}sffffl�����������������������������������������������������������������������������������������||��|�|�|||��|||x||x^x^c\^cYXWWWX\[ZW\[\\\x^^xx^|xex�xe|��^|||r�����|�����������|���|||�|^^Z^^^^^\\]\\\^\\]\\v\Z\\\\\\^\\\X\x^x|xxqx|�����������������|�||������|�|~�||xxx|^^x^ZU\^\WWWSW[W\WU]\U\x^\x^x||e��|}�����������������������ѹ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"R22.0000-.0.,-00002.2.0020.0000.0--,#####!!"""""###$,$--,-0K3RWWWZ\\x\^x|x^�||^|^^^^^^Z\\^^^^x^^^Z^\\\\[W\WWRRK22.2.0--000022.K22R2R2WWUW\\W\X\W^Z^e^^|���������������α���������������������������������������������������������������������������x�������������������������||�����������������������������|������������|�|||�}c^c\XX_XXXLSVUS_c___a`c`cffcflffffffkfflffl�����������������������������������������������������������������������������������������|}�����������|�~||~�e^^\\\\\ZWWWW\[\\^]Z^^x^^x|x|�|||||x|�r|�^|���������������������|||||^^\\^x^xx^^^^^^v\^x\xe\\\\\\\]\Z\W\xx|q~�����������������������||�����������~�~�|~|^^^\\\\ZWWWWUW\\\\\Y^\x^^|~q�����}�}��������������������ѹ��ѹѷ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������x�~��������������������������������������������������������������������||�|�}eecXcXXZXXXVXcX_X_c_dcdcddff}lflfffbf����l������������������������������������������������������������������������������������������������������~�|�|�|�|\e\\U\\\YUZ\U\\Y\\^^^x^|x||~��|~||^||���|�����������������������|||||q^|^x^xx^^^^^^\\^\^x^^\\\\U\\^Y^\x^xx�|�~����������������������������������|�~���||^^\\\W\Z\W\\\]\\\\v^e^x^^�|���������������������������Ѷѹѹ������������������������������������������������������������������������������������������������