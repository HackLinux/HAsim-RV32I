�a�I�G�d�� �O��Hg}9!n�`�/^�6�5�!q�����WP'#P�c0��OG�d��\Фs��u��wt"���=�q�8G��Si����U�/�$f� ��V�=��?�;��l2�ICŊ��/��/���ꂇ�yi�(����������<[��dؐ�(�U.q�ޒ�RF)e�"���]��/�)�ڿ�v �ɨfѰ_�Z�Q����IL�U���x�ǳ����Q�|��|>�Uxj��~��
��Y/|���$e�/����Y&��$����E{ET�rq��{��w>�\��S���,��j�O���2ȮW�#�-�:�(�6 �^D��L���y�+�(�_�\0�I�ʼ��1||�>`x���A��a��m(�Ֆ����ڑ2ڂɣ�4%\>If�|p������c�O��ES~�V�+Ow��O�{����� �`FsG&k�����;����K`�0d�-�Z���Aw������}��>��Lc��N2���جp��Ñ�|���ơ�@�֙k>���+�ߙ+o�묪�A6`qKU �!w=��W!�0,���a��9��ȫ����v��|�d����uI�܎� ��O�H��gސݯ��THL�F5�hqe��$y�7�kܭ�EM] _�G������	u�Y[i�A�lڦ䶗���P�吖���аp4/�9�}��u�)�0df\+�u��W,�� ��+ ���Z{E/m�k��S����o�-�{�X$�t�K���@)s�+�#�_�F�ׁ�
 ��n�]�vX����"�)���zͰH5����W�j
l5Rz�;I�8o��J��,25m��~�>����L6%� �[ة�yxA�GI�̻����rg3�u��������1�z/�0O�%d��Aˑ���#J��פÝ:Xwp<�����<��8������03���ŹV�q�IK�[�-�'�/�F�aW�aJc��B����P�ؓ&ٚ}�}�@f_@�ƈ��r����k��a��]����;[޽D��v�f?C�k����x��]�<�4�" 8wA�x�?�zi��?�"\&�9�.x�v��Zܡ��	oS�`y���*����5lh[��@ǐDގ�����넓�{'����}b��'��ɽX_,���q"�Y$	!��>�@4���W�)-��
�`O��ކ^Wk�� g����݂���j<`7ٱ_0����+�Uʛ*%���y��F���jxO�⬽g~����)K&�ݛ�����{�}G�A3�ϖE�(�W7L�ـ��cv���i���"7b��SJo�B�ْx��"����$�/,��Lc�e�MK2-��'<u��q5���ɤ	��Ā�ED�Q=�l;��>�=�^�	L:�I�,�[�R-��[#�B�}1SO�%Z����w�~���RǾA��7�\��U��Z��X���weBp> �,ͩ	gBeS�rN�l��+)�<�?��W�BMૡ��z)sMۑP�;���[��DQ�����x�9����'�+$`��U[=�@�	\���]TW��hR�o�����[Y�M�OJGw �G�fY��2��fF������:��`�:x�F���%'���[�D�G�8y!{�W���"&f���ȅ��^�包�t'���j�1�4x�/-�O5OȇX1��	���m�OC�����&�:��#J� �ڂ��)��>�Ue�lJE�41�Rʃ�t�&�7}�v�x�6ޘ[�pz\7���{�x�#zu�* U��pX����a/�ONdrj���Jx��N�և�>"�G�ł^�FN�yX?�l�\����`�:��ijkDԧ���"��[����@�Ď�-je׳���_�E�X4;J������@���OD����ͣ��$�V�XĹ.��okm" ���&�&�(#$�=Д�ݕ[��fG[�ܴ[��~L�T��ie���]�M��"o��?���Ye�uHS+f�@�8Q^������~�m���z'ǚ�����"&�4��rJy@���u���m�2�^m�����ȣӪ�U���}TAЛ�y�qN!�6x����t-սئ�"����*�����$FҢ��᚝o����3�s
%{����h�mM��п��F�uH��(�[��1�)ٓ��p��ݲ}^V�w��!"��~Qo'��2��Ė@��*{�\��R���I��:"�ݝ$H��`��T��̿�-d7ڄ9�y7�W��~�~]x��Yѭ^xp]�5�W��!< �}N��KP��!J��?!1O/��0Q	��O!F N��f�g��'>�`)"�ьs|����_��
�����ُ���A?�nS���!ܞk�Dڑ*O֟�wO���5���7(:�pl6(O9��z<�0$`�*5|q�R��[.7�ǃ�"���N_m?F��5�g���}w�����Q}�5��z��l˦�~�Ol��=�14�v�'���:��50��� ������"�������a�R�T$:f�عҴ�t{%i���[FF�S�la���We�4d�f{��
��}q������j ����\d�U���L����0ʟW�'��>��e�l�����7B�Z��B�WE�L�' =�]X�
��)�+Ş���0��=��XO�;���$����k�	�	;|]ʳ�[�0 � ���3^X_�F�*Ww����%����KA@��7��7^�П241��;���4=
�f�$)ԯ�t-����#�bzӆ"o�ւ��}fZ��Ɍ7���W�*=�Xc�u7�Gd�dHF��#pw�����;Q��:�+�E�3��hL��z3��݉������A%���+\.�CW�����*�nB
�4��6���S�T�W
sOD��ȴ7�52�;Q�Rӱ����E#N��6m�F��3�� �"D6c�̺F�I�i�5/����/�!<L\���2��oJT�8�.H0�u��6�*�};�k�
�ֶ�RL'��xcD�$���¡��2��F���N:����U���~&=8@ͫ�e�� Y8/No��^��{�#G,�8G,2̲������x�?lҀ��$׌55{��q���V,}���v=��!�{��/�*cXk)�Ȏ�/[G\U��U܌
�cT����~ٰv�e-�ܳUq�L�g�E�	GG���qG�W6�!����� �w�vJ�����S� ʌF��_G]�� R  si�m�  s0Q����ͨ����r'�1w�=�,mz[�!,��,�b*^%��֦I�2��%[q{�g���(ƌ* ��c/_xN�(��/�mܳ$l/�y���x����.�]=�"��
?��&C�w��pw)�V*�)��-	�zߏ��� ĞH�H���f!�k�B"�
}�1vg�vPӷ+��r;��2.:��js��Z�ҷ^�x×4�@��+-�Z��A��j��H��7�*m�5�����oGc�����0&|}�2��;�.��L�7$�(���S��� ��w�µ��&;wq����V�	��t�p�P��E�e�q��s'�ᆱ߳��
w}F�����������3�jhҠ�#qJ�t�s�92HگW@gU��{�g�☡"����j��j��E�3�ǚ^@9���˞��O5`�İ�����[适!�h��D��k�0Nzn��6G,��z.{��[���`X� E��@>���I�����e��>Blb�`������ �VH��*�D� �i�V��q^v,e�#�u��>�+�.yC��H�2�ȽJis?����t7e�q݁*�-�w�n�ݍ|"�\�&��Lh"�.����ř:F�z����4zE
�z�q�t�e�]�c+#ʧ�z�jK�j���љ���V��v)�4`a�6��t���8�J�1�z`F����������/�@��C�k���>�	���������}�^W�=�E�8MI���qP�1l8��&!_�%|��U���1{�_��k6�,�x�;T"����T�$@u�kn5'̹e+�I_-��Ҋ��j,mr
��Qd.�/U�����9�ME�.�O��+��t�z֩�J�����Î�WE���RP�䬫$�z�A&K*d9�>�f�[�8(-�VS��ҩ����o��dCd�%�h������?}�K�޾ɨ�����v³��Yԩ��Ҵ,4l��G���Q��沶��{l�K�A���b�m=pdy(��?�צ>8��7#�L����|n*�U��y���Pp���E����'��h��վ�CB�n��f� �>��il=�3�)��!S��� ��9������8?a$�Ă�"�!�wk�#l���g�VG7�!�E�k�
0�����R��}p�̣�0�����\��(m1x��[�W���#Eq��-*�]jw�t���=s[��u�q��JV��Y{X6�Y .�N���n�]�ݔ[i�o�^"w[?&ՖIx"��e�j.�eh,U�2s����c�O����W�V
|�%3h}=�W+�C�,�U�oy�7��b�f2��Y'�h�I���.WL�#|TTO{H����/y�B�um)���?q���<�Q� �)�����20�������ׇ�W�X��v�lK�{��3�7��Q���<��A��xJO �
cc�u���V C�a���ˆ�@����0���U��؁#�8��P��aiB�7�f�41;�h�$KL� ^w��@j���hiDi�G0ǈ|��w�����d��`y����&Fecq��
�<7�a�Ӫ���Z�%�����m%�#rm�0��W7�d�0�
���9�w��>x��a3^�p;ڍ;�'�J�I���Ĥ�#����e7a5�=˙Hk�c�ZLf��a!�_�/h�2I{Im�0ʐ�&�k�o��`N�1��a!�z
q���R��?X���5hY4����'����>Ǧ]D�l �9+~2,5�/M��yO��T����z�k����c�T-�оܽq�
�I
������L�)2�-t�H6�:�U& ���Li�
h��À]j�*��Ɍ8u`�|ٽyd�j6�&�D�s}_jP;| ML��QQ� RE5�D�ٍ��AD�Ĭ�8��y���l�L��V"Iݕ,��`�Nk��X�0b#�}jC�}�k���"���d��$�"�X���v��ϴ1%���
t�lz�R`�Q	�>��U�x
��8���O
wܗ3s���@�""�sk>fn6�;��n��~4����\�6@��Og���fQ��<�,�����h�Xl�R�!A������!#�z�<[۝�+BS�ѯ�Y�=����噠��������������/�%���A��,2���,T��� "7�]li_bu�؜�2ϣ�s��-�*P�+�޹mdӹ�,P�p���A�i7Q�e�jD��W���K?N܇/��>-�����Wy=�=��IN��F� 7D���J�ÙmQ�i�L��Ӵ��;�#��pl�7��.��,�'F�6��t	��9�R���0M!$O��#���*)���SR�4����T$��w2�M9�=�ǸI:>�d�!\�-�%�_׵]4�G��$��/��N ��u?�y�wdN�^>MZ'iV�m*<s
�O���{[K��������@3�3�UM�o0A���$��%A����-�I���lBx�����-�R묘�=^�[u�s�|�;0(u�p��[��G=��>�גU����KGh�%茇����;�C*(g	�'�R�V�(��ɢ�7o�Ի�������t��Rp������d��n [
���
�g����c��W�K��@���G�vk ��t�����:��"��~�oDmt�������T��
��7��2
��p�'�=Fl�3G-N���l�<a�b�V�t���?|e;P<�h-@>6��F_i�HŅ&K�T��q��4��7�՞a��ב�K�k<�)({�U��
�z8��(�.Ӝ��̝d��v�b���1�j�u��C=@%u��Q���~�����`-{ ��%�=�҂�{�N��m*�6����wa&�[ ���¬&:�F��(��i0�s9��r�>{�g�#���� ���۬�j�� �`<�`5C�>�Qr��e�A�V���?�Y��t����´�
�1��P}"��E;U���ds�ɖ<�{�כ�|��q�G�1&�v�����j({���&�Bʀ�mk��7y�������pc�S��=�!��M��k�O�+~�˟qU7wX.����;��48���YѴ�Z��}_A@z�����)�LS��љ(��@zw�Č[�r�m�*����V��q��ښ�\�}@hK��-����I����@э�#If|��3�	kvT�Wm�v�֢y��x?�u����7w�I*�b$�ڤ( ��7�h��_��	���t
+>�xm�����L0�-U�t�nC�G
���g����0��+�,�gS����3��7�j��5 ����x��B��Q��q�[�(m�?#	�Gȑ[�'2�D�a�ȅvHo��.��a��z�+�vx�55@�QG�8�{w&�yYr\i�u�`�ɒ�zbtu�W��R�w�,Hr��m.�8?�G�h'k0�7��޴Xy�V�9]����5���+�z�Q�,�Mr>���
��u�e�T�J�=|9#���dP�����F#c��Y�E�ʾ�+w�5��FC��)�3�+��`�xW��Y��nP�@�3����Sy�_�X�5��{��Lਬg�$�+M�^�	��ep^�E�nĆ:�`F�N�WClrWČt�/�i��Ic7�m2;����ǡ�����E9���V�,U	{�׆$����u��^���L�N#G��l+���g�h'cx�M�,��~3`��'��}Ú46.$���<Ϝ�|,9����L�KmSҧ>��C�z��]m��ǯ�Ռ[	y��J��e���$]h�G���Z�b{��r�&�>��VRd2:��i���I3="i�zR��y'G	zH1ʆ��g�Q��d�߲C��N�9P(�~P�`�&A��(�6��h,�a��Ye||����gZE:}Q
��k��W F�j~�|�ѳ�FS
'+Ft��I6<��Ο�)D�c�����bm�4ݾGN��>'�H�"$�go��M���C�����PZˏ69w1�Lb�4�!�	^]�Z<uE�h<z�ѢC�|S5�yBbg#��������z�ٞh_��4V�w�qo�vMs�M��W��|���3��� ����.Zꦨ�6���9O�M><�")�0�vJ���d-8z�U2�}�_�������U-Ύ�8�^��+}+$�8��K}B.z�¿�P��WZ���C.��:��~g�S�R>d@oؖ�� ~i�L���iL��$,t�em̃u.|_��-��P�}>��RP��z8;�}t �N�(HƦL��A�M|q�r����@�U�|?sA�2�1vV����E��ϝ!�ޠ�DV�F}�8�F��'�[6	�v)L��m��*�h���QOu+E��:Ek#+�v�Pzۈ�N{����i����Q0��چ��-V�Qg>�	F{�`��u:�W=�lzP�sڥ���W��$�m�N_/�D#�p'�͙K���$�u�J$e�pGl���Gʞ�n./�sJ���\��ٻr�J\KH��rx�����g2U��Un��47|�7S�:-T�O`f�:���3�V��-��ӯ�Yq�Ý\��#ר�g̮���R�)�׍�w�C}������-�uRMFXPu_}M�1b/��>�ޜD �>��D� ��ՠ>q����41���L�B4g��Sd�7�s�FQ���h_e���6�LGRJ��j��+a`]���.�����=��$*���V^�^�W��ߦ,�X��p.I�)n-΢&��F�8J��?�O��~��h!ny_Ӹ��m~%	ɜ��J[� ��y�{X\!�b��Ҋ��Yz2����i,�*v�- �B��(�>혨&/�0��d����)Dؤ~+r��.��|_���<�+!��g?��arp���=�����? �g}�4˫%��Կk�wdJ�{���Q�O�^�Y Ǽ� um	�k������qˉ+� �"h
����*N�"�a�E��;M	;��v��	Z�{ڤ�)�[�b���U��#�[��^R��a� T�b���u�L\>�$U/X��	K,d���g۟`JE�5�����T�D���5�j���D7��´��Q�c�ނ������������X}�E���H5H�fL9�n׎^Հ'�O�Ls;���"���j2��j6.����\�OW���-�ǌ���0Kݧ�v�=�(��3K���-�:jx��
��	ط%ƚU��d�@�4;Uh���\m\����&�F�ʊq��Ǔ(�x.1�d�و�N)A
Ί��{�c,�V�W���r�m;L�7/�"�߲��$��+W�묳�/$<vz+�ր�c��gF�:jA1�v�UBy<��6�Q�c�Lb�^���{�z{�e�d���^�cq7��4�c�W?��v
�&���*Vɱ��КEԋ��'&����U��1�r�����
T����Hy�=��9i/�a����;�W�1�$E�~�b�*]1L�y��5创PH�Pe�����D���G&�@��"�'Q�K6��ld,'Ik�t�&xoJɃHe���!��:�dh�������<�<����Q�Y�X�|O�E����l�g�����ą������a{N��!9�&��E�h]忓�;)_{�c�}2wD�Y	)�Xt�Q�t��($$>���9K�.dN �Ϗ^�Q�J0�[]ԋ�������6���z��RK#;�k��z�1"J���M��i��|�>dV�2d�SΦ^�i؛��Ɲ �'j�s�*�@�7����*!z/OǺ��ت����#&�&J!�>SR��Vbui����VC��܍�B{����q:�6,w���o\	��%����o��D���Vr���W�[?"O�$ ����K�2��\ʹ*g�&si�]�������J�eM�ڍ�&8>�@� &�>v�O۶%̀"9���P�������dYi�|ĖD-�u*$5��,�n&c�D*�ˆ�|
&8��?��d!������pYAw�Mx׃O�=Ľ�b�7��]?���TR��h)��^t������E1P�V����5F`�N��3P59�N�<��،L^�6#�'��(}pH��o��H��& ˞`Ic//�
��������^ϊ�%���#�b��^�� �(R�US��>9��)J���B&��]g�^>�A��r�uM^nX&�=�ctK�z���G ^k�>`�;�4��8|U�3z\��0g�B�d������!;��?K�4�E�\�lR��/е_�~6��V}~�:.!ˑt
�:��W.g�����L�M^j�v?ǚ+@���T~���s���	8��ƻs����"yc���L|:����c����3S�Fҩ=�9�1�1c��ɓE>̣��ᖫ泧�;Aś�y���_����kx!70�b���)�U�7��kS��5���2��3�Q1�X�x��R ����F�*�`#6֊�Sq���߃�����lW;�اD	5�j��Tp��.�A69�K�S�+A}-��Pk&e��P�z�������5�R�Eqho�^j��l��6���΃[���I��ƎK����!������T[_ڦ�,S�"E��Y='��CK�[�����/�*<����n3���c��p�4�r��z���J���J��Aid�q{���㢜�y�$��AUTh�B���,R�ɭ1�HF��ފJ�<�D]/�p�=r,~�'4�� ̡F��Aϴ9l���U�tdXC�]�gC4a{K&|\-�u�CY�*K<�yx�@|�����^��0��n[��q��($��L�H �~��P������:X7Hy��J�`ކS��Vt|`/9y��q��d:1���T|�I��!گ�i���Do�����|Bv��x��� �ly���pg4�d,�Ug�5��5���ݔf�ADg�*.ç��i��Wگߠ��	�����8���[f=Œ#���T�M���ks�$Ǖ��o�t�l�/��(.s�%�X~���ɳ�Q`��_b����Q��z�Y�(��۸v�m"4$r��UT�hb��/J¢;x̚Ǥ!��뺿��"W�jw���I�*l����`if���������A�a�F��ێ��H�Z��V>�p��O��I�(�7�b�ܾ�Jh=���A�Hո n����E��o�Uq�H�s�k���j�2�OJ2ȭ�2��yA���2H�)�V�ە,c�Pi��IAS4N� �O�Se�Wh��N`��H`�P	��͹�/��ѿ��K��b��,� 0�"�
�����+Ѫ�a���c@�>�Kt)�8�`y�p�9�$%�ꯤ�~"�m�\�+���O`�oKk�zQ&���곐�NQm�d��=����h��ov�W�ꝣ�	=Γ࢈�T�G���rA���7�K���bÕ�Xk��~���j(⛪&cK��u�:��-bp�#���q�Y�'��0IA����5}�5Z�X
��)�C��u��r������V!x�SG�ܺp�r��
\E����9���O������"�nV���#~�u.�`�G5��w-er�~'��E!/����m>c8L�s���պ��P�ٹ�U~�	q~�u�#�uk�1S�KT;q���Scm����)Eh����J�J������EA��Q�-�z�^2�U�6/=sm�@�q��~\9C\�����Y %~n�u+	����`P�f?��K>3�3۳Lx76-�?��O�p��UR��uW�������]%�����w����������FM�KA�T���2+�*N���U�|�4�5�Nz6�pJ��c%�U?��J�������x­#�"���#*�#-�>krm�K|W��$s��ZU��)�.���]z��Df���
Tl�A_-�$���k��1S	��ݐz\
�*��g\w�A�E��d%�����H��d�B����jp���m�\�B��z.��7>d�N.x�i"�����<����$��$�k�̺�/�2���*sewK����u�Q�_2c.|�	��I_��6)�Gp�Ez������=8�����Y��[��KT�]N�9�Ne�Pp�̤A~�s�z& ��y0E^zU���W*�>74�P��T�T���`���LPi�iDy�Q��Wo��E�}<LL��Kwqe�zO�.�χ!��`�������M69{�U��9}���Z�����<�qu�F�د�dkZ�I����]K�C'��S}p�P�~�,0e�%q��7V�O��thn�����c��:���<��1,���YTB��y܂����Tϕ�V��LT���q	6B(ޏ<��E�cq?>�tN����J��y�$oٰb���Y�fr�J)������uxD'"Ɖ���o1��4�y �al�Б4�+5� cK�V�d�C/;�j_5�����x�0KM͖i`�%u%s�����&��u��D�Yf������d��z�i��� B�ld�<��e:;��dd�#���IeB	�kG]颦��ޭ�/���a@��T����泂*\�*��#NS� ��٦�)_׋�N�>ftCx�ɣ�=W��={f�Z���r)����}��P��ʘ͔Ͳz��@���.6�`�:0����,��r�w!o� V����8�;�PT���a��4d>����[G�/q ���R7``֛$���xO��ŻCྣjJD@�x�+�@E��Dh�nS�[?�0�fT�qZ0q�I��h���r��S}w�N]�u׊7�%̏��hL2���B��ʤND�4[��7w�]���_E
�=-��[?�q0��&O9�o|��@U_
㓈.=��YW<����܍�+iaZt���F�_��q@m�ȗ-�8�c�z�<��QC�����E:��z�C����ŀ�ŉ�*��ۻ������(m��L��u�,"���t�h[b'�cY�2y
�s�����}�5�������!�mZUU����*"e�lF�Ñ���o����Iǀ����+��o���U`-<l�T8a����]�o<�0c�>WS�S��*����8�h)��ٚ˗��E�g�ct{u@$����!;Y*�cuD�r`f�����h�,av:�� �y!v	sĔc+��oĕڷX�}g�C���ig2k�tS�%e@�`�!�H ������{�ܢ��拟�F�n� ����]����	/��s�Ff���q5�a� �0�RN��g3O����Ч�� �G�"H����'�9���\�,��2���Ss�� \� 2�Ak�JR���Po�wae\�΋9�~�_&���C����h��݁ƀ$
4ʤg7^��Pg�J��^�'ۑoN'����3��PL7p�z��6a��[�]}��Z}u����eTb��ė�*��4]���W��k]I�'�b�s�N�K�بk���/[=��֩��,�9���:��/�U9��Ҳ3.")�,P��ǋ�ۅ���;���:��N9%ۡ��M�컘�i46��'3=�QR��O7���R�BT\��T���]�h�qP�l�褙HqZ��ݙ�~R�h�ob��`�|P�l��8��h���zϭ��E�{��&u�w���>tq��m�%t1V'���b �M��x5W:�)���&!#L����|��p� ��� ��#������K��J�%zF��[�U���M�Xf�^����_��1�/�p�@k�q�����rn�(�mߖã�B %�qP	��g(q��tt�C��A_�_������b�VGP��OAa��x)r��,� $�IyK�Ȣ�Q(�u��c)�a���; �\Z=��.���Q�q����
o��hI	���]��I��%V�#��9;~N���(�/n<P`�nFd��>�����	���m�Sb�JW�#u�>�)wv3y�v8�~�3peo+rwQ4�؀p�Si��v�����y.P&��+t	n�YG+MUPW�kp1V�����&x'x��x0�`���rVӎ]]ԌߢDO��68�e5���������2�c��Ďͼ�pW��-�|�2�䛕�7	К��0 �=�c2w𝻩;��e>*!7���Z�o&s���,��{)�=*r�k��+��
��4�þv[���Q��.���z�OW���_�3xk(!j�_i�3P{*�ۼ���N?:��N�I����b��|�'ե=*k��?������*{��eݐȯ3q���+Ynm�ZS�F�Gnm0�ʔ������j�
+P&gqV"���GKjFWNS���w��kn��'���x;�C�����R�\\�9���_C�8z�tg�C� �,�. V8Ȃ�J�_��J]���������|y)�ey��G/�EwN�"0�rQE��!l��U&��Q *�n���>]A�mE��Z�b�cO%��>�G��z�G�Tv0���*�BY�'16��+��슼&ȉ����,7�ڗܲk��c&��#k���\�-㶴#��&�(O:��i\�x���*���_�V�a�^g��
o��|�Q��1��ď�T0'�yUt�c����}�f�DI��bQQ���Ύ���F��4����
�T�̹-`je想re��U=�k�Z�BI���7ޗE,�������'b+���:�q�:��a��*X0��n��	2����� �5`��''ЙWP���n�!P����1�Y��׏35�OK�2�XF�g4�/ՀOa|�|CnL���t/$�s�_��?]�_+~���ւ���B��L�an�
�
V��X���^P^(~~�Ɏ�� Z8��|7���vH�f�s��U��U�$[����-�����Y$a�u9��G��l*A�z����h�\�	H�@�4�Qൠ1�a�狆h!�^��e�Q�p\���IY���dӌ8�z�A�6(h�v����^ �`�6�:=+��O�	�=�k�v���u�c�^��C�%�>��K0��[F�x�_�����A�8���tG��I�?�7��>bUM�z�1��	VT�%�S-~}�i|����}�!p�4�;���/�/��M}+]ş�y�X���S�X'Q����}8�-��6�󽋆EQ\�a��[.p���%pf]����;��U^���#;�oǂ���V�Z�T�{����´5����4��2�y�W��WBq�K�f~�$����$bּ�׌u�������v�n�c�!B�2xa��j��� ��	�I�ǃ��I��l�
Nء�7/�!��g�k�A�k���w؝Վ�|.�L���Ev�BmI��-%װb𨗆q] {�J�Cj�i��0)���<.��8��E��뜪�+��/}��(bY`;D��Y{��fT�8�S}��HD''�F���~m�Y���r'���na�M�D��o*�Ġ�o�]T��H�
�mv0�5��������g�N����v#�k���K,*
��n����T�駓��p,eZ���.������NB�[*y>����JVlJ�#X��NֳM�/�x�Lf��1�Ho��.Șr=ߵ������8}/���(�����;����~,!/ld����-l�����[�;}��9n$��p��l��<ؚ�^[��u�b�������fm,���|)�k-����"')f++�/�!/`-�z�)��!���L{	�Z[�=��c�c��#�fj������ �v���H�F4�\�"!��d��\r�����r�
�1��%ʆ�!�H�7�[��;�@[�h9"� �{�^�¸�1�����QZG,�;<+�ո1��m�G�*���GifW��t���ՃPc#�J���=�4������hi�?gtp�K>��Ѣ!.�ŵ��DU(Q�FO�Z�)��{�&e>��5��Y"BO2����V������cֵLyL��#q��_���QX��P!M�u�F.�Ә�lSqMRn�ik�9�M1cu0)�"�����F�~�q?� ".�q4�K�%���O����O���L7�mL��F���+b�����/�ؐS�}��U����xZ�z���p�ǴT��i�/U!�:1>ՙ�������
�.�4�,������Av�T��M��{gw�klқ���Zڭ5>�~3_��yQx4ʈ��u�L��x�M�DKyˈ����QP���^�2)��~�_i�+� ���R���
#%L����������,,ٳE���FF$&��f!��ţA�[z��f����q��m��l����n�(O�~c��D�����|�W�����f�V׳�oګ�<)�B#~աV��VA7����غ��vC`a�������u�����4W�\G�2�mx� +�J��V*O�Y�#>M�-i�+�ȥ�D+Vn���.ݩj���F�wm͝����d#�	ӨQgE3U��_CpX�aȐD�yxtY���&�>�E|�CI*D&.�2����p��{I�!���ꈌr�9�D� �"mXW�0`E{��UC���Td9kDh�I�q�\�����rX�)ԉHD~s�5�vK�F��VweOQ�v1Q��d�|s��!7!��?k��P���v�l�Y�csXW��&�H�}�L@��8d����zW�q��ɊE�)�8����o{` �SzUh��ZU�2N����r$cf�s��c䇡lEv[_W��9�%e,>n��
��p������U���'��*�Ѽ��0���������wW_{uP����u4WTa��p�5��}��$�yr�v���1cJ�o}���j-�8W�Y�s�2�U#9grw�b!�R����,H�i{i�b:�(�=�f�D����ՉN�>"��or|-��圪�$P�8��}D���Ǜo�[��P�@,%�c,Ya�"m����#<�_�����sxC�amy_LPk�b8=�4�oulԉ��e$�y����2��+O	<u:3X:�*���������4���0&j�vW�XԨ>%P�Y�{��~�x�@0�Ҕ(Qě֣ā����T�Nc��c��wӌ �>GSf\N���膟�?em�&���-�I���F�Twx���{~�4)e�3��'إ��-�s��Xg����x�/
謯�w^p��g��H*`+R;���)��!���;.����VP�-�t cvzh��ѫ�\*���� k�5eA��ظ���>��;=�Z�ڎ$�?�O�7|~F<ef���&�v��Rz	�3��~�f=�p�34l��6}�.e�)'p�N9o]\äBz���� �Zx*L��+����Ub��&u�Ŷ	gh.��L�4M:����H4�Ő�t�P�.-��� ����+��%p���cB����vO �Y��D[�R��=5��5�q�c�E~-{B��"�ٍ˜e�|-O��u�+��'}�8�N��з}t9`�Ǥ3&��^-�G�ҏX�Ƚ{v�����C�����>���UP�FK��fE�e��Z0@��"�h��c/˱6���2Ӷ5��e������ i�7���|�T�+e:�'*�:�?d��˹g�~�m~;��Tx"⃁gW3<#*�M�cm�4���ݵ�'(t!g��r��6����×sԒĉN-p䃁��1NlMb��ږ�%�O�����au�e���X��'($��y~�ʳɞ��D���E���_���Xο�t����X���x�tk�$u0�t���8Gti��pE �#�;��p����1 h���ۮ���!��	�����Z9ȑM�����'�f��������Z�k���=�S�!靱��J�׾���7R��{�UU��PU
�/X�6�¦�S����
�_NNU��ȑ���%+�|�������H@�Ѹ>��P��F�ɰ:�f��^&�c)��'�s�xVvbخ�ڙ�1���!�뒗k�N�HJ����c��6�o���f{�����ބ�=���o��D�1=l���!�0V)������@o��TW��e�0�r1)M,�j�-*D~
6?\=��|�E�Ю��5�\L�'��0����2�G�!6���k� ��S���~�u����[�������� U���O���c ��Xd�+��j�Ur�TP�u��R��%,bK��#uBTd�i�M��Ke���W�rn����ĸ�ЄQ���+��F�g��K퇋���Q���c�U�1; �����u���kQ[�tQ��2=⭂$U��.���=�]�t6��o/��O�#&�#訄x��N�l���6�.����z���i�� �^쫳�k���P���v���_