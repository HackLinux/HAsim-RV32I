���������������������������������������������������������������������������������������������x||���|~����|�����������������������������������������������������������}^|e|}|}c^eXcZ_ccXcX_cccdccdcddcddf}�����l�s�����������������������������������������������������������������������������������������������������������|||^|x|�|e^^\^\\^^\\]^\^|^^^^x|^^^xe��������������������������������������|�|��^x|^x|q^^\^^^^U^[^^^^^^^\\^xx||xx||���������������������������������������~exx|||~^^^\\\\^^\Y\\^^ex^^e|x|e||��������������������������Ѷ̶�̹Ӹ�Ѷ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������x||���||����||����������������������������������������������������������}|e||}e}^c^c\c\cXXc_cdcffc`fcfddeff��������������������������������������������������������������������������������������������������������������������~�|x|x�||^^^^\\\x\\\\^x^|x^^|x~ex||����������������������������������������~�|xx|^�x�|x^e^^^^\\\^^|^x^^xx^x�^x|������������������������������������������||^|q�||^^\^\[\^\\\v^^^|xx|||�|||���������������������Ѷ���Ѷ��̶�ѹ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������