��*��vw��R�;�2 c���q�����<�Ù�F��-%^�le�=�dY��E��z�T9��3"*���%jA2U�eg�̨�ԧT�^q;>z�_i1�B�%�6�T�F�vV�p����f��T1�Y����!�Q
��\7p]���gGmbC���g��-�@V�����$�}^�?���Hh�=U�%uB�H��a������ߨ���E�ŷ�pA�`�TE��tE��f�u�/%Y��n}�@�N}� ���!猏�p�_`�>�HQɯ@<�6�)O��>�,QY!M��S�c��䕎0o���\����<�%�at����=�"��:�J��j���������#C�/���#d:����B�dA���!{�eS�[[ ��0(G�RpfjG�ݐ�yw��:bQ�d���]@Է�C@Z/n\�����m��5Aeb�C�AcE籁�å� {������A� 2��Ls�� 	��d� ��ƭ��#�KtU.��r�L���^��N�����?g�pd �a�}����:���Ώ^�ΐ~Z,r�n2���O�������=�@+��=��n� �M����!�@��뒳=I`��N�<�!x ʈ@�H3���i��m�2(# dS�/n�_X��t�;S���qֵ�&�l��
�tayet���e�d����MH���X���r�b��J�֔�)����JK8fk�2x�d�k1J��@�n�o���
�{l\㈥��ȟ��G��ҜI��O�q�w���)"���-s\rzW�+=P������G:�^�_��_�ݾ&���_nXf�*$�z�g��b�Е����@͈�B;3^�������)�t�����^�x��&G@�-K?�:�9~�qi�uR���er�%�[��F�Kg�HF}�N&
ws��g�6��xe�9�*��@g��/�1]CD{�MK�����@��g�ʯ���aA�H� �©�- �z�e����}��D�H��Z�zYA�����̼F�;����C�NT�˼�Pˀ뫳t^�5&#�9Y������+ Ƣ�T\M�8�{�t��/h jH��)$�y+O�K�7�{�Uy"�c���)�K�������
��j���:��f$�[@j�k����L�;ũ��#M�Z}5d΢�Q�4[O�A[��,�=�m���Q�K�� ����%����칧�؜�^ڬ����r/��0��D�j|�����
왆�A<��} q$hy�������]�F�� j�L9�V�${��R�W΀8�!���Į;V�3�K:i��|@�����B��F�p��w����.����U�g��������P�Z�'�lع���M��B�����G�V}~@5��6<��db���&�G?q��ˊ-�vg0��#��Swhh��R���,�3�l������Zb�m���b{�e���xhr��h����e$��[dҜ��[�0B��#�����������>���ql���(��%&�|_H](�B�͙6u*-�cΏ�/�l�rؠ^#��Isf��!�)
�
�iש L�D���~:P���u�k�p���.�i�J$�K��허��X�tp��^z���Ǧ݌�.�W���yՃ�*a�H�s(WMI��wP��_�(��Tt|j�Dy�;��9I�{P�Ѡ�򯖡�ڳl�&7�H�i���4Ym_�WH�]���P�
�轾�Ⅰ�f?a��̑���/��;W ?��m�i��9y�H���?�jG�Di����� >��G*�?Wo���z2�g3,��PB���U�Eu�'pr9V�3��dBYf��Ru� j��4�K����%s�9P�b>pE��ڿ��d�k�nsཀྵ����H:W�i�/�3W@�����]���_���m����3�2S�#d�b�U���$:7�=�@CX���#	��&*�
�S@�5�h�����3e��f�l�~��e]pe5�T>��J'"�&#.3���%��������I� g�SPwW�%�¥8~bL�L�j
��s�C ����%�oZ/fU���u�xbzi��Õ�{�a�����"����{�e�&� ��w��H>�4y�x%H��k#T�j�瞽l#W�H�w��mwR<'� =��U�|����]Cgg�=�X���AU�:x�&���LVx�T4�늡����׋�z��/kt�k���|� x�"����*����2kY�nY�QlYuB�t��iY�c�O�z���s�z��_fǗ��`O�����&R�ˣ�V�]�ƎA�<���Kdګ�V�D��}���V�|R�rU�ĳ��e���a ��&�ֳ}ě�c�e4;�b�B�!�)��v�����ɣ R�A���l���g��g%x�R{����0��74ȋgEt�*Ng�)z�V��9&�3Sp��?�?��Z��R"#R�`�ԟ#�|���=��T��#�-~�Ը���<"/���o ��oY蚍l$�0ם�/S�*�X���ou%�9�`(Ď)���L�d���0����$Ԛ�v�f8�'���S2�_�D���-�h�7#ɧq#��b����'���M�L�|� �K����R���Hj�`&��Se�M�e��)��d�#����=,���n?��܄��]`l������?��;�ek�����z�b(�b�R���s/��������;�mHn�&%kSnqSn��یNnQJ���E�#u@Rs�]~�7���M�%y��.S�#�P�ӟ�����*�$��Y$ "�ޔ��ArE��@9��f����4Yԫ=rz���dC(B�Jq;Jr�W�U8�a�����<��עS�$�Xc��IpS�N���G�n����}�����
��V�y�^^16���	����4]-�;g}�$����xу!1���τ0�)�=�Z��A`lsY�ň�w�]��d#��<�蚌�w0���EZ`���fi�;̖�ak�$ɻ��0����XP��:�!��������_�zb\�#��Yp�6sb�8�n����>��9e�8�}��r��k��]$������R�� hi��hϛEH�-L��Dߍ�S#M����}�M'����ϭ���>"J�S�B��{���A|�׬UԬ���5�PS�����'�_RU�m����z�h�o��գ��Y|�%���V�zvs8}��tu�� o�f��d�N�ISwsh��$� KF �*�g$ɝZ6X進��X���OV�S[J�����X��giS+���g(-WXV��IB�\$�u�;Y�K2�eQi-�,a���8�Kk���ݭ')�n(���#�	z�dT.���B������Ͱ��D��5�}��=3�a+������a0�N'�?��n�2����cOJM����B�]��-�4?j�DK,z(>ұ�I��l�W�4�s�6�.I�w�Y	����Y���u���ظUq6XɔPR	,3�(%f
��~�+C��;j�*j�ϖ+�((FդQ�<ϣ2�SȔ���U1�Ձ]PlV�+g���A{z?W��H;m��<x9���&:@֨v��c�W�-��v�H�������M*~��u��s�?�^=�諰#�o ���-O�{�,^�Hd��J7C
|!Nt�$º���p��^�ԙ�4�MAj���Zw�b4:�@�A_�6�L��-�Q=�~�В~���T�T8��B�$D�	e�UNfFM9�4����ܤ�C�����4�r09��������>Q½�+	����;R��G� ۝��D�}���^������5>~�K.E�
!~ͱ��p,��~�ZR����E5��>	�@�7�fd�_p��[�(h�_G���?7ܘ��{���m<�AF�|�0����t�օ��=�Sv�{�S1�;�]�w�P��*k��1u��`Ex\w��.I�h{�,�N���EvX�xa�2!RB!�K�ji�{��UMh,"��gv�Ё��w;���b�8F��!���ʁ��,�5�L��Wu2M~�E �sV�T�4ָ.��6�ɵh�z�R3������H���e�K�jT��0����Z!�Z�[4�Ԡu���N8y�)Zl�ب�c����"[�_q�E_�0o�^_jo��Y�K.��.�(?�B�d�`��I߹�QF�|�I�s�vq�/Hdd/���$�~�)�3�E���x�1��g�{ ��2Z���_���k�Io��_�����1��Vb�����R��U��l�d�F�}���'%�6���#�e��"d�����:���읧�
&Efӑ���!�_�6\
�"A��^r���e�X̫^��r����*�G�G(Ɠ��j	�vaƋ���� r<�w!�*t"���/� {~mƐ���c�X �E�x��뛓���뛓�bۿ�����`����`�"0�P��(k��_0>��瀖�Oo�T_�Prs;����}{��Bc�z����dbPr�|�pO�z�f��-�z�� ����_�on�E����wΑ\�p��6�q���i �Se��������#=e�����v.�d,'��� ���T,'���Bzؔ@2"G�'.*#���ǖ!�^b�����ԛ���t&�j�':�&�[nꛏ��C������ �3kd��ѝ��<cy&�p"&�Ⱥ��a���[D�����Kb�Ku&�'n����B�&��#?lל`8�s���'�>*@"�h�B��`>̦�mf���E���}��z��.���u�BpR-3��պ��� �q�m��a���ם� ��ղ V�(]��'��\�f�}��>� !��o��g+�5D����ꛣ�&����	뜲�c��:mP�b�D��dS����࣍�)���e��*!������Ű�������I%/S�͔<�i���d�3����Js'�H����d��q �����>� !�<^_�ӻ���N�s�b���T�*i�*��c ���뜂�c��p'�H $�뛧pb�C�b��t��oZ���b�C�����c^�cޜ���D�V#c��X����&露�c������ed�5��T��%��G�d����e�-b��-���m0ǐd>�>�^��5��������b�f�/9µ�����"