$�~����?�c2�mT�Х�%\nB�Ȝ���LR8G�+�GQ*zű���,iQ7�R�nO{O\K���S'�-M����Թ�;ow�J>tz��HX�{��{����ɸ1�aL���Y�5 �����Lf�9X����|�)�kJp�������i��fV%m��ڕ��2B��`���%V��u���~�DhX��I�d���}�X��)#�n8���u��)
/��Wf�\O��z�����o�g��z�>u�zb���4y�E�=���3s���@�扡+�����_t�Ql�e���uC!�+�Z�+KK���0������]�K8�t��:�c���i�ΙC��s�������~\IW]�ѕ&]m��gP3��'z U����ӵ�3�ub��p�^���#���A�ߌ4��i��I������8����_���GG�Ѕ���/�3��0zqrqf�|�-0���:R`�FLm��7q��ZC���6���m���@� �]�y�|~��:���-��ʘ}[i�W�7�>pq �����'^N��A�}ۼ����<�#�;Dɫ,�*�(��"�CC���/{��x��2l
��C�x����
ßn*�O�o�_:��G�1�?��8,�A�k�)����� �;�&�\?tl�X���s]L,��9~v9p2zm����^V��0������u���j�'~}A9<|"�E�ډ3߆{�x��7�yt7w��a�$IW.�kolbKGM��ޠ5�Tn���?�"=�ͯ�!�
�ٱ�U����k��·��앷�x��5e\�˝O���h���P�vl���L)��\_+�5�h�kf��"���["�]�L�}�\Kx����ѫ��/�u�������Oii4�4�n�r;Wg̀��t��z�O[�Ho�	����i^�է����J�(=��F P��p�L�8���>L���R_t	��Ut�.����ȓ����O���8#6S9cW.`�h"$���WM�.�7ƱU���􅨘
��_'�W��jQG>̦����:�%��ע�"�!zƯg���wڼ�m�7��-w�7<O�F���(7�U.1����%��L1�B��R��%4�#J�������@����@ˤ���bK웚��#U�5z;�1����}���'�l̎)Sz�PA�B ��{�M5Gg~�����Բ��2�=V%��v�.�;���0a��������"_>��p��~e66������m�����Y�f��b������t�g�&%���4h�z}h�=e��(�3� ziX�����wO�I���wO�Q�q<�d�D���c���x��&3��4�:�!�\k�V+F^kU&�m/<ް[���~랦!ؼ5�Y��nk���'�Ǖ������_����"7��!�X�Ӓc*�������>6��x��y����݄�$��$�P�9$f���bF�Rƌ�3�&�뉌�&��-V�h1%,-�<R&�2eQ���� ��"�3��HA������Xp�i�`���O��X0X�%� ���C'��@�ā8�;�������{���HŁ�o�8J�st��Xy	�8��b��
Ҁ��/vO�no�2��)
.Hc<�L�e���s�����^�Q���k:t`�K�1^^������K���4�r�m�����I��5��pM�nl!�"�	E���+-�4J	}ָ���qC�p#t�gT>�cJZL�M���0��B��1���*��8�~f͊f�"Li�Z�\m]�k��2�:�<߱*���K;2���XS�!���O�ȼ�Ұ���'�>�B6�:U���l�٧{�RC���VY�;K���<�Q�OWp��.��zT��N7����(v�(���
�~M�ʙ}qL��f�X��Q�Z�rZ�!��n��x�i㝖��vǷ�_bѓ7���I(��D�&FA�L��ur����f�d�Du8ڣK_8�GT��vP�E�cǾ�m*Ș&N�(]&����|�#��e���T�X;6��(�ED/JL�u3�.ՠ�D���ř�45=�(����������a��-,�w�Rƈ%sG�E'+�P��O?���C��PQE���	�}g���=��J{�����{����O�G�}?N�o����OA_g?��&�wl���ێ/�o�Eq���K����	���8�/�٪\��;�n���}��{~�w�������9߲��0pw�ć�b�O�K���s�]_*�^�yo?�-x�a�k��4���R�v��[�a��y���xkl�1}����g�o_|�[q��E�������|�ُ���Wv�C�� jNawK�}��?ʔ�Ta�S�u�g	t}.`��#��{O��׬H��ԣgD��ό�%��p�xF�%qt��d�k*��n����xY�E�Ⱥ��8��i|?d��{G��U鯑�6߂�짴�+.Y.QT�f{�re�BȓC���R����E�����h�t���>��2],�K�D��L��l+�����H���G�%�P͔`�Vۙ��JIK���\%u��P���R��!� �������Q�+@��Sa?����γ�q����)��9��o���)L�25+�ߖ��.Rѷ0R[4�1.��q��y�	�{C��T��߰��Ëᵦ6�j�-<����jhZ������Ej`;�I�2�/��G�"�:ʉ�.��R]ix1�l3��^EԊ#U,���+��v�!�Ry�^/�� �@��� �� @^�T��%����ite�Vѩ�[R��:LM���C)�_V�����}�Ϯ�I�i��Om�L��3�I��Yp[fU�ke6u��ԡzh�m~h5z�D5��-ȭ\���*x �CӠx/Ʊ�K��,޻<y��P�x0�}_3����3JՓg��^Փ��(O�x��~��c�F�2%�
DC�H��e��� L��f��B�'���ʖ�lZY�ZF�2I]���&�e�x�� ��(��]Yx�������6�Y�\<&�F�o�y+n*�m���h������n�<fYBw&�ı��a��/������J����4K�ZBi4of�o�T�WCZ�D�͕��Z�ୁE.��B���L���^�uڄ_P���%T%-��h�%$h��e�a����fj�
�e݋Nt�	u�$�b�_�&��b�b����Ju�U\@I>Q��*�Xz(�'B����51��1��= �o�pW�ڌ�Ã� �"�:�'�
��L�b�nIg��p��*d��r�����G���⼱�A���GT.�e��Z��!6�^.���z�g�����ێ���u.���"]o5��\�k��Z��!����q����-�(�|\���yT<���	��z,��lM0�˞��Z3P �.����=tm�iqkRG�|[o]�
h�
mrA�����y���=uv~%�J�6��|e�	���|�xz8�ê�O+S�� 7U@�V�g!?�]V-���>��~��Ps_���+Vu�?p�"n"�-<��mL-[��(,�+����s��%�:Ǣ�aq���5�6�ldl`R�}f�j�>���D��aOr��Sz�cL���O99�3'�ᰜ��s(i�M�F;��,,���Hc;���D=���d9�/0�����8�TX��
}�r��������0�x�6��kd]Q��i^+�g�:��۵ǯ��D4��7��d!z�'@��]i+eoDx1��~�����U\��SD/{��e�qR��g��
���JP��Z��\o�2JfL  �&��
o�ZO�6bw�̉46�+�W��׫�#ͨF��ڸ#Q>X�6���2��ޫ������g�Ǟ����`[�X%�S�� z�'��Ӹ��G����H�~b4���/(���gE"�F�קoڗ���atY�w�~B��0��;��o�ٛ)��|����.\BYŮEV�Lp=1��.��P�U�����&]�yf�<�Ɠ�f�&��>'�,�8�ӯ�?�دnd{�v V˽��h�VU�/l�HK���P'�z�<A�
�u�n�����6řx�D�jYm����2D� �śL9��e�~��ņ_US�BK>PK����xY�rӁ��~X�f����+���^E�����ڂR�e��(���jU)�yy ��S�%��)�
/ߔx�T�`9;[�_���=j�r�*ި@�VpH�I�yR���ǣg?��J�q�q�X��+�	_��~[v��ym�g۔]�cB���B5�~��g�E9Ҥ�gl���-ɱ�3d��|��Vq����Xg>����d�Red	}�a�����<���Tfet�+�apDɬq�΁����)������e�HE�to��pk�?h
��-q$�����-�Y�"�_L��Q���?Qx��z�2��R��:_���zz��ⱚPl���;C�7��jnm�y��Z<�Z8��8��T��c��W�YV�4�c];?�;�hs��
�u8~!�.tC���X��ʭP;��]U�a�</�>��ҵ��CC�3��p7-pl�R�m��)��U�1�7狓��M���`�:��!�`^ud~_y0�jZ�GW����.]>tr�ۈ�"#HR�)�V���V�Tw7%"�ʲ;ۯM/<2ˈt�bL='ϧ-���$"1�7%`��rc� ��RQ�S�#㋣C4w;=Of��AG%6K��=�q8����!".2��>uxָ��zEi�H`���O���y��Dy�MO�Lq��)h.��#(���Sj	�O<�kn��V�G�鉙��}gŴ�J=��2�yc�0�����1��x��&�<?F�_uU+<���2K���L���Xcox���a0��y��ًm���#�K%�_~�����g�R��]��ư�o��}�r�Z���F��u1�ψ����ϙ���n�&q�s �O�о�=�4�7Ƭ�ZUɉ���T��������L�BC�҆uW"�_0=h��Ics�l-�|�7џ���
G|
,l~�>f�W.���0��.����}�x��4� �����4mU>���S³6����e��gϛ.�F�b�i-�?
��H����,�Wi��K��	+�r�q�'M��u4��LA;�D��E�R��$|�ګk;|2��[{t�mC(Y�2G��3ONd�zū[{�4�>���Jo����{�P8rC�1u~��H��NX)�^>;��U��A������z�R��!�������6�~���1Ӛ�ȽQ�,H)�Q\{����F��Sh�?pWB��5�I�+���?�5����4s�1w�
?}A���)]v�轈5X����OL�&��ޗ��ӋH�=�ޞG�ɼ�kL�'|G�I)��#m��'�(W����~��]=�F����i����5���{WM�ղ|���{����4$l<)�ݕ��������FǇ���w}U����{�瞪8|4�W��ًiv��x�R��2^�Y�<h�ۆ���!�|�tyq��/h9��Uޝ�2�Ҫ�ps�_�_�t�Ce�Ǎg:��5���n�!�C�������Y	�4��4H��ZL{?:��Yq�֧�i��.Y����*�;�Mk�2)N�~��6�Ҳ��9�6,����-p�0VԝS�������i4١�1���A�Ju�fu�Z=�a^�p�D��`nq��n�+�/�|��O��'6�eg�D������<��\gJ�Z�Q�s�����{�+V��Cl]d��r?D��eU2�/}��Ե7�����>Jk�AֆV��Y����H��\�Q�Gj�1������)�#�p�cfս����2i6��7�ㆄ�퍿�*7��7����
�4vs����:Ž9򤢳Q�����w|H@ˀ��,��ǒ��̀��@��'�WuC�Q�a�bg���U\�@#�s9ǫ��~�\S�����Tck��!J���k�Ь���Ep��
��p|C�#��4�Ad/��V�h�� �L �Ї-��� �:F �CK�}|S��ڦm�@�R�B��Uq���(I�ҚRH@l����s(�BٚZU�.������馎�/{�o�Q7��:
�)B7�u��ӥ�eVZ$r��9�&i)n��&�����w���T�ڦ/�'n�9�����$0�Q���V+�1�ذ�zhw�#��
Q\��9n���p�O�C>}iFh�`����S��4瀑�]L:�f���'E�q����'5��ҵ�sH>��`o��h=s�49���zd�1��d�O��r-�N�O�~����X;��X�63j�l9i��܃Z��sZ{�����÷��߶v���6��ͻ@k��]k�&>Hu��]���g���M6��<RX��#����fB,0l�%<ʹw�>��C`�o����.����}���s�j�Zj?ݟ��E��<�rJ?����L6�Ik2y�.����^=x��v����5]/��J3�I����j�����y|)�v�>�jC��� B���5���lb�t��ԗ���?-g�7�8l��γ�_�.d_i�r��[����C z �h����|9`$q�l��p�aJ@�?���B��'L	��%��j�]���XaO�ќ�	@h�^ۥ�>+��pBz���2��GH����>���i��.a�݂0����aܧHNgi�"���L;��X0BIU��ԥI��e@�(Kd�mANqkR����@�='��F�T�f#Z��4�fһ��ͤ^�7v�6A���m�gT�fѿ���W���Ζ�JK����"�X���w�Z �/�#�*W�f�V��B��a����]��A�Zm�NϘ�B��^s	���<G��3!~�oH��6Z�g�Ǎ�p��Om�o���0�,o�Hx�MJ:��s���ۘ�|g@,�ʋ���y�$��E�*�j�2)�l��o��.ޮ��!�Lytђ�����}�D��ވa����.��?9�ml=�����ך���ښ�:-->ŵ��gܥB����|�^:��`iZ�a\���z	�A������N�}��1╉Fq)���8�q_/�6�Qi�V�Ԫ�x�y�L�6�t6���!/-���ҵZ4<����Ϊzb�n����N��[�m�fu������*�m�Q�����'萲4�8�����e���L��X�0#ʞ��E�%��4�@�:^�(�/f�rΈeij��м�B��VރBn�P)c���h�= x��F��k
L���a6N��r�ă${\�b?����U��nz 渦k���k��5�i5S�v��gd����VZm�ݢ�!^����9k=G�k_�𣷐�&m5�E�q�rtSw6S=�����&f�R���u�/���"ɽzy�Vfg��}pC�`�z���$2��u[��yE����I}��3dRڊ��T:��ipe��\�_�,.s�\�&M>�+�F�Ɇ�l��O7���۔���2�
V���sߍ�e�k�ڑ�Ȣ݇���/V��١�7,��� M�(<�1�^dd��L�P�\\�8�O7�L{�>[7,��M>���^:�n0���0l���އ��!�;W�_�Q�˃:�� a�]��ڔ�S��$dj%�(����PaYRc�S:�e�z�}�>x�]~�5�L�bi��3vJ���hn��-�&��^B=��1�\�9�Q֎
�h�:�J-7�ʹ�"{�F˅����ˉ�ͺO�{$��.��b�$:�Ꝅ�s�n��?p�Y�A�ԫKV'��hɵ��	o��!Ko'A��t_�pm;���Ρ�o�����<�Vf�B�����-80������=�ie;"Q�@��A	���Y���䚜z�P�N~~-�Rϯeo1ne�i�S�ݬ��T�!���ϭWԛ��4:�ք߅����:�w�0�z7 �e�M��y���b�{K�0c[˗W��Y*+��$��m6�t�~���8�]D+�)�eHw@�	9�%��ؤ��AS���XI��ck��/~N�?T��[/X}٠��R��������?\�)�y��ـ��\�.=��qI�3�{��ӈ;`5�e��7� ��	w�$����qpK�������f��Ӫ�$bZ��,C]��'}�fVU P?. ��D�Ѹ��ۤ+m�#�E�$%nS�.$lf�drꀨ�%�e@�� �ɲ7<zY�9ҳ(����d�l�$51~�0?���/�D�H+k�F���ղ��"�W�g�w,���m䬐h��������h�K�}H���S�5���Π��=<_���'q�q�h?����5)�o�R ���%��@�I8#�S?(��C�HzM�B��&��w�_�C&郤U���|�@d܄<m7iȯ�#����]T{x��% 5$i�1n���|]�/�l,P�*�x�A�M*K��I�,-�c8?v������PUU�8�Q�`M�e����wD��
>z�Uw�6C���}�%.���7]r���Z|H5���.:�3fY�����]��Q�OSL�u�])���]$kDkf�H���dk�? ��yn@�&qx&M���L0�#Z����2�����T�[����B��_ئV]`\-'�Ӝ�+^�	��g�D(�V28(�k��;������%V�ҙ�2]6�1}@I����/�����M=��v`������OG�<������r�&�������G[I��;.��LCן:��.��?�#M?��3<��p����i�!11��BdoE>���X~(�D��8C������X���ߧ
�mA-��q�2V����<�}9q���\�E��]њiU�A�~(,� R%��ϑ�yu�M��D�>�R��GQ���P�C�,�TR�&��ōU��������YF�"�H^Ԯ�����~�^��W'�����������f*jP׸�y�i�=�~y�n�K��[�&h5 ���%r��V��*-�37�I4����Zb�|��jK���:�Q�˥�}o���Ey�sq�k�<4�Y�6gY���k��?�����O�n��6��i�E��n��l��O�y��Լ���+���
�b�սA�^���fc��Ƚ3p�2J�;#L���<�(k}�:���A���p��� M�$u�t ���'m�T�UK
%��`@.�����!��<%�u!��;���zV�=���m��Gpv�x���R�f�b*��+�L@����=(bfO^o�F���joK�v�Yꃭ	�hИـ�3��m���c&:ɿ37Y�K�����3�3��i�����)��g̼�,�8��uVyKb\"j�qp{W��qqJc���������7��)��6 �����
�H�7'h���l�qdd M�4u��������W�_���KkMe����{	�x���"yy1#�e!vO���4�P�%Ugb�m�VS�Ք��N�a7�2��f����X0ߡ�\P�l�I��:Us�}_;N��r��F��)1�/`�!��b!��'��g���i�4�p!��M,�V���w�Ą#ş� jF#TL9� h�]�����i,�/hy��ɘ����B��+�DO�(G#�=F}�RM=U�J��7Z��_W���'؁�0:���(:�����=-rt��I\����'�iX#):]L��Ϙ����L$�]���;jMh��������?���[���ig\W ^����ޫgU&��ؗ����9c�����Z��^i��C�7��C��u���U?��j���Gs���<R���=1{de�-��%���Z�#��J\+_O*y�WPO
:&���yk�E�}�s0����\������!m�I��/>�0�ع�(������{ nK4��Ϳ��Zu�x{�ͶJb)?`D���mWi�mZ��߾4ˆ��v��Hy�]���O4�����й��i�_�ړ��)�~ z���ZI����Ɩ���CJ�x�
�B�:I����Sf|����ͳ}�q�ݽ;�M�u#�N}4�qO����p� ��DV͐��E��"���?f���a�b 07�V���ijg�2�6�U��'Q-����`w��;��)�U�p��?��,�� .��O}=D�0���̪�i��	�I|�,7sB�YZ�l^(��䓞m	�z�+�>��F��K�5� �����UM�&`w�O�|p� {�:�%mR��� �:��.p����3��
m>
�8@'��3�`�j`��w�����Z���"MKlj�V�$T���I�l(z��Y�	�Ԏ8-�!AM���O�t^���A>l� �hu�>�VkO
qD�3�e���q�[Uo�[0��Ӥ��A��..�	T��1ŏ����H�ѳ�,��Ʋ4�����[.D%tTIV�r��|_9K�l��U�b�RbZ�t}F�42/�4'���ig���	�gy�}~�L$M�Vʒ1�sC�W�K��V,?��m]�$��"���zY.�WU*��ȗ�n¬
ЦD�byzv���Ɣ�C���{���h$����"���N���6�t�$�Y~"������	����KLI6��l�tnz�*��8䡧,��fDڐ�La_5�)�cw57�ڔ�i��p/H�Nl�j$<N���5Y-�dQ˭XϒmIQ~�_�������K<����?	e`���(�L?z���X��ӫ���c#��X�X�4��33�`T��2s��m���?"ŋ=�A"IDý��Չ��nn b���q��n5�8W��2�z�e���}�$&�{���8�Ί%�Qө{��_�ōDI�v�Z�i"5�:��rUdocP�w��^��Ỹs���s@~�bA��ᯚDV-��9�ό��1 ���[%17�Z���g7m�U����yx���ޑ�_��)aR��%o�F"{�>"�Җ"3�)0S�6<�jVӱLe(}�\��+E�k#��J��ӏ���j��bdy�M���oi��PR}X
�~� ����3��ܡϷ\X�.m�[]jY����twlm�y��Dt�G!�X�Tq"�S\ۨ"����9��1v����[�V����p�4<YAj�'�����{&I�뒾�cj�M��H�͌mp��18���ɽ�����Z���.�e�8y6Kl�>s;����i�x�8�mo�,�8F�EU�-��ȉc �	�����)�Vt�N���;]y�<�]�b��^�p�T�M��gWU��<Yui�`�SO��t>��O�b��銸ѺiѤ�v��K\����_���6Vcm��s⢆jhm�hmj̵9(�A{��~����� �M�����ɕH��,�@.�ro��x�.�����{���a�VT'V�K��|�;��<QIS����ȍ-�:	��F�5���*����RF�[*Z6��OI?���;�>�\^⹌�pR�%�&VGu�����
�~�Tmj�	��=��m��S5�&�@��E���ۂ�('�V�� �E�P{��2���q����l��ɱ��'|������i����|�:��*�E|(	�X}�L^�����u�;��^���L2��β5a��F���\K�ޘ�)ğ����B�_�u� ��{��\�wgfuFN��� lz�v�$�s(�2��|>�V
�^�1$�?ܟB+�w�p@�%lk�o�~�:���&���Mq�� �s RO��e�F��1�+'���W$沩�O��P���!8�ˤ�x( �܂=G"̭3Y�����j֧��Q��B~+5�nV�u�4�r����A�<z�Tfݒ	G{K[�D��ݻN3wO~q@
7�]�Pdo2g�O���s�+r�!��^�+��Q<wH�Ы�:�	TM��2�9#X�_UR"mn�=zo��������G:jQJ��{k�hc?�Z���8U*B�6ڣ"s"�c���jͩC�|�1$u�| F#�.̾[!��F�]�jv}�x�}ܡ�����Yq���>=�kD�0��+�!��=������4��*C��Hx����,Y�e���eG�n���	4�k�2է�n���5�A���,�p4n����uޗG��Rgi&cPċ��i���6|b��»�u�͠�����3��A3�렜�z��1mU)�v�E�����v���K��1�!���KL�o�!9�)3��<���)^��f�:��a����r��h��}w�e?���m��v<.�Hޫ�6���}�D�� >-�a�qV	$.�S��;��]L�n���C�$�9LS�c�}c�'�^�a] ���ZwI-S��lJec,�R�8ߦD]�}�*�?*�ZnUU���!v�x�A��XPؾ�R��}�M�$�]��7<�ܰ�z�d�45P� !N���K@8S�;b��y.懿��[q����k"?~���Fz�ad���#ȉ�Xr����`��f��+pG��;]�p��X�6�ޅD�o��=o������@�1h��C"��
<M����w�Q�m,�4~�S��qd�BtxdEA�-v5}�n*@�L��+K��ss�*~�ܹ~g�X
#Cx�H �-�b (D��m�2�)s�4GG	'���5b'���zT;Z�S-�J����lN.ė�HW�0�V����b"�3qGy�BpT���a��εoЪ����B˃����21Jc�xS]-�'�zw�,<o�	�#aUi�Z�d�'�6��� fP�_*�A�x��I�FC�-'f�ɿ3h�<�+���fʻ���[6�gYL�Y�>N'�}i��Ӆ�^'!W�Y$s��'3;g"{�9�SU�q8_�ո�d���9�$\v\:=#X:����g����7rrCG*���ʸ�l1�fr/�~��$"�r%��XZ��K"�4��)>�0��x�(v��;3:��W��U6&�� ��u�Z���!�r&�Vi�Ѫ��W�*�|��y�eோ�{�(��6a�Hl6r�H��}�o W����Ef�v$B+�t�㎺u���z t,��o@?�@e�ye̢x��E�L�k�y��w!Es剄\B���23)��z��;Ƹ1?Y�6��M�h�*(����|�W@�K���DvV�VJҵ[+us��T�ex*�k�>��__>˓p\5�ZR�`H�T��q�/�)�������r���-��.k|v7��Ε>�`<Ns�k=#���Ie�[K3��CH�H]��ڙV&�i���vB܎���-+��~����M�v�"QՇ�)Ώ�h�}|���+ q�#�G���m �gc*�Sk���Fޒ�/���b�Tg�oiN�$i��z�����)ה�6�6q���8jv�ƃ�����+��V�DD��%m�Vc׳��u�������4��L��P2#b�ZT\cW� �@��#�Y���m{4�]�ӝA�Л*��O��ɇ�G�e疁*c~��Q5J�1�)�\�\�bo��!�Pk�wdaot��j��r�g)Lf��kpT��p/=�1�Ż�kY����9�gKh��6ǽ��x������{w!jX�R��ƚFY�=�o�����.~	�|:N�����E�+Z���.�'� ���'���n�.����s���h�� ��]��-�o�wm�(��T�ۮ�Đ4�XD^D$�Q���g��THB��Sw�6��D>���B�}m�e}�bD���M��c1�t�9��vm?�S]�D�����nE]���#�y����>�^X4w���D�"~�fE�����զd��wJb�zX�{3���f�nˇ��%95�5��[b�E�¦w*��Eo��}���?�=`,]�G�4v>Otލ3�ۧg��0�Ļ�� qA���ݗ��=��<�ݞ����<�W�ݞ��
��7��)4}�R�fM9&a�mq���g6� sw����w��� '�l$j���/�Vi���$hᓜɳS��X &���m��Q�#Z�Q9�/+q��3��0B4B��`��U� �/)pm�!�)abW�4&����J
������5��;iA�Wˉ8������&��������'��&�$�I�t��������$�4�30�ƭ��^�f�����p5#�Yר���ʅ�Hx8	��g��I��}�H7-}��nA����̃�����W�}	r_P
4�YI��X�P2h�fؼ���`�
��_�q�<�)�x:X�'>	�� R��	#�N��2}�_�����wDW��s��;���v�~	q/��3O�qH�Y�����e�v�!�s�^��'��bG��ڵ?>+��n>�'�ƽ��d<8�<���}�x�b��'Y��[������/�h��8"�8�o�C�9:?��&+��8���V}�����Y�����y��R?�[�{�Q�Lc�&�v����X ����`@lő�\�J�v�����d��(�ltO�]��%��~����mҪ��m�з�� �ʠM�:Vi�,׮���q�|�Eoz�;��a�)�o����D���K�
Tf�%*T2��@�kc8��2c�S���c� 2�X�pEFo$遖�؄(���CX��Z+������u�Wz�1S�yF��Th����u�*��v-�168h�:3ZN�S3���Kiz��?0��l�9��i��yH�J