R[9?]~�ɷ���P��භ�ȶ�Q�W�|�|����A����B��\��[�^������ߠ������{B:<�YyO�U|��[`G�Q��|Bw���X��y\�Z���ߡ���d�����~W��~ݘ�z�o�uªm<��W���R}tMt�VtMV��tp�pppJLoLo�oo�s��q�wq�wg�_��WY:8[~ �4�4��;���4��ݘ��Tѭ�l�r��y�z��z��f����چ �RNZ:9�~^^��A�Q��E��X�B�śQ�[~�ƛ|���A�P�yy�`��Y�D��z�����������{<��Ù��W��[��E�W�wyWy�yP�y��_��G�����G�ׂ����V:\@�T��TN�umm�mosp���c}ttVtM���M�vS�tpM��o�LoLolU��qwWkw`Uj�\�\|9Z8[~ ����ܒ�ܬ��3�����T��r�l�ݓs����u��N;���f竄��{R989]~�^W^��[^��\���Q�|Q|Ś�\�^���Q����[�U�\\��Z�^������ߢ�����C����ǚU�����E��^���|�ȖwZ߶��2ָ�Gק��FG�d��ˤ��vZ:\|��z���s�<��u�sq���R}Svtt���M�Stqp�t~ёN�LLools��w���w�U�jBZ�_W9ZYP~ ��4�����4ܩ��r��J�T�TT��ܑ��z�ѐh��ݭ���燩3��lR�YZY]Q||������ZQ��ys���ɟ�]�ɷɛ��|����[\�����������8�N��ނ�����C9X��XY\�ęyxA�G�~���������\ȵ���\�G�eGH,��F̂�����vA�8�~���z��Wu��uuosqk��R{Mtt�V��q�pqpS�Vpё��o�oLls����Wqwjwyj�����w:Z8[~ ���4ܒ;��;43�r��TT�ъr��f�Nu������?T�hhff����; fR[9Z?�ƷQQ`�[��A�Bs���ɍy|wŖq|�|A��Q��[[y�\�[��Zu�ʁߞ�����������{9u
�?Ҹy:�U�``�^������[|V\^�:����GG�GeG�d�IF�Gˤ��V~9:~T�z���wm�ux�osq�U�RSptV�pqpp�qpp�v������N���k��W��gWwj�yjw�\_�y*Z8[~ ��ܒ��44�3�������TT��J���L���������r��hh1�fګ3� �CC�Z89�����[��B��\�y�y�B����Q�Q���|�W�>���X\�O�[��ʛNǴ_�Ƞ���˜��� PC�<���E�Z����ʧE^�W~|��ɔ����``��6�G�G�GG�de,�b�I�˻�x{�::~��l��o�Z��u<�sw���R}vpttjqqqppSjqVt~�o����o�zs��w�jg�kWjUB�q[_��X:X[~ �������3�f3f���T���TJ����T��zzo���TN����������� �}R98Y�W��^������E_Z�úʍB�ŷ��^��Q��]^�ɺO�B�\Z�y�_���N�Yߜ�������r }}98�c�X\�Z���QP��]W||~WV����^Z�����eG�eG�G����H��F̠,���{Z8�~�����o�Ou<��oswU��R{tSt�jppjjjqVVMV}�o�o����l�p���Wq�k�gj�\�U�\��X�P~ �h������4��1��z����T���l�l�u�zNoz�zzz�;ffګ1����;� mR�89�W���[����^�֔��[Ȗ��^�[���^|ŷ�]Q��|��ZZ�\�y��ʟ�ʥԜ����칬���R~9���ԸP�XP��\�E�E�W~��|B~��^��߼7HGeeG���)�eed�d˹bbb��{B�@���z��w��usuusp���R}tvtj~jj}~Mt�t�}V�L��No��l�}qjwkwjpqU�k��w�\__>?E~ �����f��3㬬��z���T��J���Lvsѐ��LNѐ��h�3ݩ��f����� �R�Y�PW������[�^�����\Ú���P��WȡWP�~�Q^��|�B�Zʵ�W�Y�-�������F���r� CPN��-��/\���/�^]��|�|�ɶ���Z`��H��׃����eed�����b�̂��@\VT��l�Nwx�u�<�s���kR}vttVVg�}����M�}��ooo�ouo�U}Wg�t�gjwqwij�>w�\[߰\~ ������4�;3���LT�J��T���h���{��yz�X�����h�;;�㫫f;�� �C9�[ȶw�[ȶ[���\�[���=�X��Q�^\^Ț�ɷ���\B��\�A����ʷ�ޑ���������;���Cuc��\Z�Z[Q[����VW�}s�����֡�GG������F�eFe���,�̂��bI���Q~�ѓz���xs�usu��w���VtStM�����jVt�tVV�ou������wt�qj�w�wj�w�jj�wj�AߖP~ ��1f���4�3ff��������������t��t��N�ݓ��h�������� C�~|�|�^�[�^���\ZʺO�ɡ`ȶ����\���^�[���[Pߛ]�Z|��]���D��bb����՗� CNc���PP������^AV~~��}����7�`���H���Hdd���,I�I����������8P~�lzz�N|�xOu�w�WkR}pvtpM��pV�Mtp~}��o�om�No�spwwqgjpqjjq�pjj�qq\��E~ ����﬩�3�ff��zT������ѭ3��tL�U��z����h�r�;�����3����C9�[Ś[���\��0��[ʡ��\��^�\������[[ɟ��E�[\�|ŷ��Ś�_]��������������CN��Bȷ�P��Q]�^��V�VX���YE^_�̓�HHe��d�,ddI��̂��db��؂�P~���z�N|�xyx�u�V��U}pttV}pj��}}MVvVM��o�o��ozjvVp�p�jjwjjqAp�j�q>X�E~ 11ff4�44�f3ګ�������ѐ����w����N?��z�ݐh �h������ ��� CYQ�ȶ�����ʛ�`����7\�y�P��E����^͡�Ρ��^E��E[�ȷ|��:ʠ��������՗�4 Cu�\��\�[��ɟ͟]VV��V�~]��ߥH��G����e�)e��,�bII��I�⤗��DP~���z�N�Xssyuu��Ww�vVtVvq��VpVV�~VvV���om�uNLsvpj��pqjqqpjqq�jq��q�2V��f�ff1f�f3�f��������ѐTz��Y�U����T��?ݭ���㫫������� C9~|P�PP�[����[�\�����E࣡���7����[����_^^E��P�Z����D����������4�;�<�y���P�[|�]H�]�v�}}Wƙ�^_]��7�H�e�dHe�e��d�I��Ib�����\A~Jl�z��wx����o>V�W�CVtM}pp}ptvVVVtVv}��o�ooool�t�p��jpjjwjqjww�jky�g7V�3���f��3�f�f�����T��ѐr�T�}V�Uz�z�������h�r����3���� C�ƛ�A���ɷ�`���[ȧ�B����__�^^Ⱥ����R����^���ɚԵ��Zǵ�z���̻r������{Nc�^���P��[�͡]�vVV������\��7�Ⴣ�,�F�e�bb��Ib̃�IbI��:PV���z��|<�Os�N�V�W�CVtVpVtpt�MvVVpt]���o���o�l�t�ppMjjkjjkqjps�Ukk�j2V�f�fکff�3�ff��l�T�T�Tю��LW�tuW��|�ݓf�zګh���3���;�� C9~|[�W���|�[���ʸ����ʸP\�Z�`֣�Z�H��ॡ�[��[��X|�޴����������Հ�}����]����|�Q�]�}~{Z}}|]��ɡ`��΃���eFeI�d�eb��˿�b����P@��z�T�|xs�U�NyV��sRVMtVvvvtSVtVVV�~�o�o�oooljtqpp�p�jjwMjjkqjs��gs`V f��fff3�ff�f�lTTT�����z�я�����ё����瓘�fr�f���;��� C9ɛ�P[Q��[�Ⱥ�P�ʟ�Y`\����ֺ��7�������H���\�\ʞ�^�ǂD����̠�⤗��u�O������|��^��}�V}�]]�}�ͼ�H�����eI�,�b�bb��I�⹿�:Q|��z�T�wO��x�?��@��R}ptvt}StSt�vttVv���o�o�ol�tpqjM�jjjgp~�ggk�skkg7@�3�f�f�f�3��r�ݘ�TT���ѓ�T�{MuU|�z���z�1r��������穩��CY~�P������P�`�`�ʼ߸ȸ2���`���7��߼7ּ`֡�֡�`E���[Dzޠ���b�������}��w�A���|��^�]|vV�~Vɷ]���]�ͼ̓�e��de������I��b��I����A|��lz�o|m�mx�uyV�W��}pttvvStSStMVt~}���o�o�o�ljtpppp�pgjSjg�^skgkK�g7V f�ffff�f㩬1����T�������r��ҴTu~Ĵ�z���ݓfh�T;�f���3��CYɷ�P�Q����P`��P���Z��_��7ߧ��7�_�֧��༡��`�\�ʁ�zD���F���I��bՀ}��Uw|�A|��ơ��W�t~~�]�^�������̓d��,�d&�����eI�e����#\A|�������Om�Xs���|���V�pVvvntjtttptt~~�L��o�o�l�Sqpp�qjjkjjsggWUMwwUK7V �f��ff����㫇��T�T�����T�Ǒ}{�UY������z��1r����;f�� �C9�|Q�^�P���ɧ�E����2��7��7��7���H��ͼ�7H���H��ʢ֦�_�ޠ�����I�����~���w|�W|�|^�_~��t~~}}�]���ɡͼ�H��G�
�d��,,d�dbd,�b�b��AA���z�osmx?xy�sWōsR}t�ttvvqnS�}vMp}]���o�m�ml�npppqMSkkpjgjkgg�kk�q`V fکfک3�f3�f�rѭ����T�����}�}]Y�z��yT쐘�rh;�;�f��f���C9}��Q�^���[�^�\�ԧ`�����֧7��H�H�HH��༧�����_���ʴ�Ǡ���F���̻���VN���wWWWW�^^�~V�}�~]�����������
���F,ddd�,IF,�d��IbZA@�ѓzToUmm��xo�}yŖR~t~tSvvtSSSSv]S�V��ooooo�lkSpppqSqgjkkqkjkgkkk��7M ff�ff��f3��f�h������T���f�}?�tuz�T����zzz����ڭr��h���C9ɷ�^��B�E\�_�`��7ߡ�֧�H�H���H��H�H�H��`ߣ�D������ޠ�פ��bFb��~��ww