c�7CI! �\�轥h;������_\�����y��<^ �+OB��G,K�"(ֽ���̊��`B�f Y��ޔ3��˼�
Ȁ��;��
 �9s��`3��ܪc����;�.�h��&`��#<Cdkf6��@�N]ڋ��Ud0�	9;�_8b�iO<f�0|v꺤!?v�Db�T0E��p<�FaD53�2�7Yλ՞�A����0#G���z�ūGC�� ~~�(��K�*�Ea������&"Ԃ5P X�W�@�� <�-��#.�-M٪� ��E]�G�zJzBv����6�?��!�W�rԘ1�e���Wi��X�iC"���/����>�Oq3 D2b[Z����T���W��
0�1�R,�%���P���&����"o.��7��2@~o,��O���X}g�43Fs�
��9Ym��&h|~�%�� P�e׃�@Ҧq�>s�e�����s�w�J)j�0a�4��)l�)�på�z�V�jM �Ĭ�s��)��Ҹ2��&1��P�������#���r���0!z7��(eR)����\�����Ox�[��p�d�P�L���UƖ x�E��g�&�O��[h9�C 	�����2���iB��	Hh����B�����ۨ��|6�yh�/4&��[;�(�cy�����V��/��F�!�������-o�x�}��Ϗ��W��&��(ty@���v��μ�� �z�i[�U4 U���� ˔�7��C���ۻi��v��m�w2b���N����v��|#\y����}%�����ɘ%�,����t֜�0?`/�'Oo0m�����Iq�"
�d2�蟲���P��y�z���V�iU�T��D\;�}��6O�nq�n�ˠ����9�!s4Wa�m�$!����7����%�V�^�el!vթ<ѳ;�z|^�	�S����!vtw�7�W$9��g�:j�f��-��1�����_�Y�p�Q�C"��	1��q�"̥Z0#� �������Xꞕ 2��2��62��/�3 7B��4+����ؖ4p� �;K�ҹ2�ޡ�Z�Y�Ĩ�@��u�?�P�.c��Rʳ:JD�U�}DEXC,�X���\z��w ��;��{�/
6���*���ŎvI�Ѓ\3����`&�Ѧ����C�&5��4s��*���_�����&������- #"Ѻ��_�Ci=ǹK�1�ݤ�7L��F�k}p4G�=}w5��B��Xp���jrBi�%�e'�z%��p;�y3���X�d*ϙn�/�K�E��׎�����]Y��TO	�W��� �[e ED���u�����<�qe�"��8�WmCh���Ah�~���+<BEi:���(�vc�$i��� I�߯h������CB��B0�4�$
�hF4 �J	f+UI��9?�A?H�Fe���R)[
c|Ƶ��k��ߏ�y�*�	[v?W������l/��_���*Z/^��@E�����5��twz��4�JO&�lϗyM��>���Y�����b���� Hy	V~l�=Zߑ$�<��_��(��Aj<��b��ªܗ�hW�%�Xq�Ƽ�'�@M�ʽ�.�؅�sW.�%�95�����7���O|�v����P��U��Ѯ�{�l6`uo=q�tƖI~
r=��	X<�m�h1�(��Ҹd���A�|�Lp�5a$ ��+�!L̺��:Y�|t�n��p�N�m_�_+5��T�YW$�π4�]4��#h���R�
��4!S�,r��31]�8z\jgL����դ<�q�U��y��I��=x�����A��o��؂��S�ٚm
2��P�m�j%T_��6�ρ<8Z�K):n�X�����Y�(PҪy-���0~�k�b���
�t�G��:>��|GV�ý��p���������Ba��:zD��vQ��0��]���'�}���f���D��ڧ8�����W�A�!���Ϝ�a�?]x�ql�����djr�+��~m����86`�Em��x/����P�V=e�n<��m��f�r�V:�aUHO�"o�xDt�yk�N�wpq>-*R�}�@��l&�	nÑ��� �%��l�.���S����94�^��i������y������2K@���G}$;��p�`�c�(%�?Q�9wf
���ȯ���_y1�l3�~�ꠉ�P_��~HBG������Q�T:���]:˵����1���qTN6m�ۤ�����쩔^*�	v�5�X!4y4s@���Z=�`Żؔ�s���Yo�����aƷ�b(S���tb��U[,ǈ���Ƀ��x��,i�VZ�;T�X�-��لݿ�:�!`��#d7 ˕�LX�n�0 ���U��QH��'nތ��º�C:�o���@�MK��t�ۢ�%i�g�������/� R2��MW��%�@FBJJ���FL��� H1��u�������'Q�����ǁ��'Z�V�if\�yj%�\�8�Tҡ-{F2�9P���I���I��4-Z� v���9�=�D*0��3g
�GJw �t�0�`��ѻϴ�>1��3�@�bK� 4��e:;i��>��oA�0��3�]  ���OccF��3b1z̹	��5IM�Nio4u�E�U%pij��i�{(�2�@�b7�����@�����0X���rp~�3�Ds�dF��\�