)���k�r�8�Ґ�eE�N�gA���N1T<P�������J~�ҹY\�G_�&�|o��3}�;���R�욂^��G��A�>A)�gqI$��0��fa.�>� ��^U�1�mZ1W��F^�7ځG�S�?>���j^F����c-���ư�&�TdD�����U�U
7�[��nh�Lw!�Io�7ś��h��O����:�]�����T���1mA@�����C�z��S��|�����^coFʈ��t�+�&�2&�����퇤z c6�|���M�#=�~x�u_�P�7t��T��G'�RSҼ�ö���rz��`�XE���e�5�T�O�9o����F�Q��`��V��@7/ ]dval."�p�˒��e���j?��ȼu�cL�xZ������)õ��IK�:�)E��<���@n������K����|{�������~_��x���ѐU���;Af�j���w��B��b�����}��,k�C�� �O`9VMk=*5a��r/\靝�)�Tp�;����tg]�D#x���I S��2\�K-K�r���;�,)R�6uN�?d��{uA��7]鑙��V����Sd�:���O�g��-���z0�A�A���h���b��s�]R���=�YY^V��dX���@.�ȯ���Sc��s�.I�ja�R�����\Ϲ���{Kag��gdU�k�͑�ك�=�!�rV�܏;g��p��N|�p�#<}���$[�r�\-w�+�QZ�C:[�����ߙ��"�Wr�]��nz��eT�s0�^�\��9��T���"��.m����:�_į�V�$M~�R ����QR�.��Ec�$(O4�@�YD^�w��hm��_�}����1�k��Ӝh.��~2SZ�
VKk,2�p�k8��u��j�!N1�:�f�SK����(b����}�n�v�m/�;G����z��ǡw2�:��}�ӃgR�����8r:��BZZ
�|A۰��I��"�Q#�-a��\¬`v�SԲ�X��v!1LGm��������g�U)�R�qo�O����C��^4P������?	_����K2�Jxw:��E?�_�aeX5�]���`5�H���k$���G�AJ�^���9p�;x�Q+g�c:Ȍ����3�����}����7��R�k=�#�m�T�%�)����0z�oQ�E]`,36ی�V�������(��tVzx�^��pe$8z���n�z�����9t?PN�u�Z��w-0�3�|��k���X����MD71F�@&J�t���q��z�nau�3�������z�.�)�꩒���̞����˵��׍S�k	�Ҡ���$�F�������h�~.�ȁ<�P��o.;�I0tc6�98�:��J����Q֌ou��r�\/���������*���	ҫ�5�:@/.xO��z���C�T���D�`u�X:�n��h:V��e��'֕旸ٍ���"� �kF��K�O�dtUW5F�SO�tK�;ܟz��̏�*��bR]f����0r�,��g��L�	9�)�)	�9*b��Lt9����|fr�����.�l����3`��HHYAvۜGN(dK5E�Q��nw�7Q����SG�}��%���I��<E��}Oc@���7�B�~*b9Q�Ӎ�n��_Z���j��R�Q�7p�u��kx��z���������w�w�;�eҝ��1�k�=>j��T��)+�K���$�HgcD���<��%��"�Ql���(�kʝm�1�5�#'��v[ǐi�؝m��,tV;G�`1e|�Y�=��,[ڭ����{m�tU��9�Ig	��]��kc��$'}�f���P�@uhK����1KC�8v�}d?Y�����C�uf^���V��u���vO�z$��H���8�+��`5R�)\T���z��5U}1"���r�:��M�����g ��+F��O�#����̤c�e��g�59���U��'G2m%���b��!���F&�����j�n�4�?�HPs����v��j5���w��r�L��������s�I�v�{���3^��˫k��n�~&?8K��?П���?����B��A2R$�y���i�����|;�Ɵ�\��(����+���8ld2]��۪o��R�%��]��p{�]�i
N�D��e)x�|��fy�D!��SUAԃ����bx�u\]C��Rߐbs��� |�>����@j̀��<��;�m��
��|��J��W�����?�^S�쌃Y��9lK�=�#�9��'�ɉ�Q��I!�����o�A�m>7cZ�,a5�['��R�9���h��&N7$���'	4���	��.c�ک^j�᥊��r������9�}��{l�d�p�ݺ	���?��<�{�
3Cy�������S���^�7��9��/-�����k��M�</�+�Y���L�������1^Y]�������j���_E~�w
V�'��w:7�P�)r��Ż)�K/�*c<f$��/�[�� ��#^T���{�� �����~E�:���J���'��.�f#�q��E�V
w�9��D��)��I��0��g��g`�Cl���o���X���v-����~bgw�w������d��'2w{uV=PY�ڻ���H��Y(ݑ��[u��(�H��'\�:|�d���OĢ�i]ڙC��I�Vl%[�α�| �q��(*��Qb3z1�QШf�6�ӌy��Fts������zI����>�k~o��:���Nc��������������|t��L�7<�__e��UR�j���TZ7�[ĭ��q�"y^U��7�[���>N嫥#"S��ꓪd�CN�44mNӳ4������4��	�G��%���`�53��lhN77�6�Zխn��k��