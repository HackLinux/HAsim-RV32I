��������ȘȲ�����ț���������������������������������������������������������no8d`W;;;q�nqa;8aq�����q���rr�ɲڲ��������Ğ��������wwwqqqeeaa^amedaYdYeadYW;;;>;:;;nrnq^88^n�����q���qr���ʲ�������ȟ��������xwwv8d2`m;XdX;;aaan^Ya8WWaagaaaq����۞������ڟ�nn��x���ğ��qqq�qgxqnbbdeaqqdY:a`Y1Xd;;d;;;aaal>;W2W;aagYYag����Ϙ������ڞ�mmxx����Ĳ^a8....;^...88^888675/...58;;88>1.8>.22^88785..ddddegdYdgeqgdgqdgq�qddY;;;;;WYYaaYX;WddegdddYegqgeggqeq��ddaY;1[



















e;gWYaYaa^^amebaa;^aaad^;;88888881;;;W;;WYYaaa^^^aeeaa^Wabada;gd8danrqq��������r�qxnnaYeqnYbabaaa`^nbd^bnrqqq��������rrqxnada�r8qaenn���Ȳ����Ĳ�rrr�rnxrqanldlnaabdnolqner��Ȳ���ɰĲ�r�x�e�x^baqhq�����������Ϟ�����q�raddama^;;;^^aqhq���Ğ����ɲ�Ʋ���r��>a8aeadYbeeq�ʟ���ɰ�gYaeaabdY[WW`;41188;YYYaaeag��ɲ��ʲ��dY�e8a8;aaWaWWWaeaenam�rggr�grgqndYW;^Y^W;;1<>^WW^W`aadaeaaq�qgq�Ș^Y8a67...18<225WWW^2;YaY[ddYafdaaeb\^;Wa4<).8a81.8>WXW8;Y[��;eaqnda^b^88>Wa8ann>888;;4;aY;XX;aWWbaeddek^>W^98;aY^8mak88/>da/a8;W;aqana^W>`dY88YaW715)811889W^WW^;8;dn__^^;>Ye87;a^^2a;a^albWenanrrna>588a^^971.122;883;24^Wbd^a`>aaibnnda8858n^^<Y/W;;WW`;;^annrrou>a_kbba`X4>488WW^YY24Q;WY;<877>ilor�vmWa^bl`q^2d;ddkadgdnqkknnmrqxxoebk^81;4W448WW;Y[YYeea`Ydalb=loerxqqnna�n/d^Wad��ro�rr��ò�qxvyn^aa`>a>WY;4a^^^abWWah��dwqqxyð��rxoxa�l8da[qndmnrqhneaaedennxrnb;aX;d;W^W4X;Yde[g\edemmmaaa^aeeqonxn�d.aandnqpwqqrqqqxw���xdnrqqnmYXYW;922YYYqmhh\grdpqmmdunq���ode�r>;W^a;^q�w����q��reaenenneqdd`aa;2WY+12;>nYWYgr����edxrqbbobd�r^YWY;ka;`amkWWn���ư���Ğ��rrw�qnnbWaW4X;^abW4Wgk>7Wln�ڞ�����n^Wamd>5:>8era^>8<8W8W^^^lalk^>>>>^6=;1)2Yka;*Y;;mm>5556299_na8n;aea>klm`k>^;k8;^W8988nll^8887^aanlblaaXaW^le4aa;8>>582W6//ro>n;^[Yqxwaqdn�qgq��ri^k8><^k^^aaX;;;^kbab^;Yrnnmpeqqemqq�^>>Wd^.aaonqeqexmqpqqvnaa^bnWW829W988;aa^7a^lboxn\eexnnreqnna>;`a`8a8�kleb��q�Y��Y4eqn�xxr�onojvooxndng���xrxngg�g��xannj^nm�qwwq�u<qe������g�����������y�xxweb^baYYax�rnqw����������������Ğx�n�r>a1qdaaeq���q�������������İsr;�mnqdX;W`meeYehbeqgr������������ugaYYYqddƯ';;neWaa�s8bb9ԱQWY��oa)Gra4T4G'dqe/yU2;WXabqa^^�a>a;;;^qqmq�O-pd�Y���eb��پey��~v׾a����UrQ�r���gq�q�x�xk�a;q^ennr�r�����I�ɦ�������n9��a��eag�rn��eq������ľ���ʲ�Ĳx���r8qe�q�����������ɾ������W���n��brg�on��q����姞Ĺ嘘����������i�nw����r������ɿ���xrb����Ӟ��r����w��q��㟞����r�������yxڲmeewq�����T�Ȳ����Sah滹nW�ee��4eS�rYU�g����]�ala�������������a;>a;;Yeq���hs�ښ�������������������sn��yr�����O�ϲ�������Ϟleaen>842o����������ݲ����r�xnn�xoornlnnegebXQ����������ʲ�Ʋ��nd;dabnqnqemWd������ȟqrqnuqqxxneaddYW4;YWX[��4a>��������Șr۲b�Wpqndrq;1;aYX;;dgggn�r�r�w��nxrrqq�rq;SY[[f����{XXYa��rqr���qaWW`YWWYae442Ya[XYXR3;W;Q8;88;;addeWXYe;444RR[xnY;4YYge[dY;;gb8YWeW`342X_da4^eqgY]RXX[W2;>>^aamaWY;24[e44***,RZdddXqhgggXaarW.Y;Yeedqdq����gaa;Yqg[dYYYY;a`a```aY44YY[\[Y[[dg����gkYY\�q\Y�e2dYer��fdqer�roa^lqe]�ffdenrea>knm`ane[egg�gfY[[[��qqaaqq���g�rWgYodenqrq��x�xroenlaYSRXa;WWYa>kkmnpqenqedeeege��q��rqnqnee[�g2nanrr��q�g����x��xunadggpmnnnnnn>iumkunno�x���ef��ǟ����qggeȚ;eaqnq���ɲ�����ʲq���q[[eZaalnnnemimmkbxq����ȟ�g����͞�������QaWfqdgegggefq������ĞqnggfZ[[ak2o;<;^``bqghgeg[[Y[�������ȘgȚYa8;W>;;bnanqqnbkq��rdakdm]YRW;S��YW^;;::;^^WWaaYdg[[Zd���qf[��Qa2^881;..8ae^>mYlaaqqqdYe`[[-ְ�addYW;W1<7<92.1;aX44RRZXa��h��Qe;anY;2;W24.<8.>an>78>Xd;a1��d��dnneda;ak>;;998Y..;XZ[11;S��4Y;W_aYdaneYa;aa^77;;<>=7_�n1*�1;8;;;Y^^>^;aaln_aW;XW1**47:>[Ya;^WYe\[aaedaX87.5^kk<76�v887�;15;WY^bnj;^^Y\Wano_W41*XX>:d4^;aaaWdYaeabqqn^677<8^Uo�1W;:W;YYbaaia>a^^^bono^2)2**X1Y8>aaWXW;ananedaaai^^^�񾾹��(714W`YXRQ^Wa>;;;XllllebY4W44;1fX)nalmcqqqq�grnx������{nan�񼮾�*:4RW`dgggeb[qmmqpxxrð��rqgge�f1d>aqq�xxxrrrooegqqnmn^W;8x򿹾O.33R[dd[d[rrg�qmqpnqoorgee[dR�;)eadbapmnreea[YWaeqrnaem;a1;��-8133[gqde\fegddm`Xdaanee\aSa�f1Yanrqd�°���ndrqqnenkddeWYa;>��2110,Rfb�ren�����qdqxroeYeYS�g4YW;8;Yaa^^^Yo���ɲr�rrneneYak>v�a;3113d;;WYYWa;;a����ʰ��r\�\W;8WWk;88Yq^a[8aa^v^aanrbYa^W^a;8l>><1001;b<4;4eY>;;;`^ujWY[e�d2n8;qbaa8>>a;^89W;6..678b^ld^>877;>k`kX11amea8;4b;`78<<8..2/2gY1n;aaYqqnqwnuk`d;2e^^7W58;85..2;..17:a`^X>Xarnnqpqa>`:7>ak68W^an>enoorra^;;nmlnbaaalkW^<aaW;81;;73<`k>`ZaZqqn^;;Wmaam>d>n^8e>/qaonlrne������xram;88X>887i^aaa8^aamkmnquaXgdg�����roa>k858^dWqqr������Ϟ��Ğ����İ���wnunwrrnexxxwqw�q����������������x�o=fW�������������������������Ę�Ĳ�������������������������������j;:222W^a89WWWakon�ƞnanluka>^^i^^^^^`a>::77>i8.7;;;^neq��wkikkl=;..).221.8.)..))/822/8);.bqqqqrrnnnadWWaYaaWeqqrrrreoegaer�����ϲ���rqqnadn�������ʲ��n8aabe���ĘgghgYaY4;^Ybeq������ea;888WWaa;YYY[dd\bed<29W;^dWWf[;^aaned8Xa7.)213WWbaXmbbd\8abY.;^XYnnxurrnd;4W;Y4S\aXaooyrrr�bYnqohr����reddYWXae[h�q�rx����aaam����������de4Q4Yn\g���x��r�r2a;:>be�qg�x��qnbW42eSSYdaqes�r;Ymmdkddr^Wkl^aadnedYndg\ddeWea.lnr�hqbqqrrallnqh�r����r�omqq�^dqr��������հy�q�gq����������۰;;qw�Sge��gӻr�y�r�ʤg��hgg�r�a.eq���������Ŀh�x���λ�������x.n���q��㕘�ַ��h�������ִ����۲a;Wn�������������r֘֘��������.`nnk;Ydf�������r��[\]������ֶ��W;4;a2^[X3X4;;ameY\YRR[g[\��[gWYqfpr�e>d]d[dd`mdeg��g���q\���e.be�����ruaXcaenmu��s����ǲ����gdm��������neZ[qe`mm���ȓ����ȸ�2878aekmqqkkZR��[Y;;abad][f����;a4a47;;>7>7jx�[adamadnb;3RR;][;WYYdda.7>;j5d14Xealgbroa*,RX*^cdagnqqnnnֿ�-3XZ]edmf����g]�Xanwxgeaeqda8wֹ13Z�]�����r��]�Raadwne��rqqbY>ư703f[g����ʚ��g2b;;k>8;<8aba97<>>03dXZ[XaaWY�Y^brnakmWa^88;11.>`XZ�qfdfdpbbW.nr�����Ğnqkkle^nuw������ȟ�w�_Xgr���������Ğqxqopp�����������v      
! $$( ((3(00!49!A! A&I( A!A(9!9(A!A(I!9!!A!!A(!I!!A((Q( I(I(Q(Q0 Y0 Q0U0Y0I(Q(Q0Y(Y0I(!I0!Q!!Q(!Q0!Y(!Y0!I((I0(Q((Q0(Q9(Y((Y0(Q00Q90Y00Q99Y9 c9 j9 jA Y9`9j9c=jAjAjIrA rArArIrIjAY9!c0!c9!jA!rI!rQ!Y9(c0(c9(j0(j9(jA(r9(Y90YA0c00c90cA0j00j90jA0r90rA0rI0Y99YA9c99cA9j99jA9jI9r99rA9rI9rQ9cIAjAAjIArAArIArQAjQIrIIrQIjQQjYQrQQ{A {I �I {I�I�Q�Q{A{I{F{Q{I!�I�I�Q�Q{I({90{A0{I0�A0�I0�I0{A9{I9�A9�I9�I9�I9{AA{IA�IA�Q�U�Y�YT$�T&�Y!�`&�Y�Y�Q(�Y$�c�c!�c!�j!{QA{Y9�QA�Y0�Y9�Q0�Q9�Y4�Q9�c(�j(�c6�j0�j9�j(�p4rYI{II�II{TL�QI�QQ�YI�IA�QA�QI�YI�IA�QA�QI�YA�YIrYQ{YQ�YQ�cA�cQ�YQ�fH�jQ~]Y�cY�YQ�cQg^�gYjc�rl�QA�UF�YI�iF�YQ�hQ�n_�rp�YN�iQ�hY�pd�gU�pa�mY�p_�}K��Q��a��q��Q��h��iɅj��}�����}��������}���ã�  seat_r               (   (  (@ (P �fg���̘gfg����pgaW5dgeX54X]XQ4QQXd�fX[[XX[55ZV]���gXWWX[egg����������������������e<4<d��ǚggpf�g[[[Wg]gf[[XXX`XXdd]egf\fg�����ǲ��gg��p������e<55Xd[Xfgg���̗ggg����pgaW5dgeX54X]XQ4QQXd�fX[[XX[55ZV]���gXWWX[egg����������������������e<4<d��ǚggpf�g[[[Wg]gf�<592395aVWa^Xa395<9<X<92+3/4<555<Xgeggpg��pgp������q���ɲɚ����ge<//VXV232<Ydamqamgp�q�medmgeagp<83///*2/92323/32232/3Wa<aXa<V<Waeaa<XaX9<XXeaWaVW<3WV<593295a<Xa^Xa395<9<X<92+3/4<555<Xgeggpg��pgp������q���ɲɚ����ge<//VXV232<Ydamqamgp�q�medmgeagp<83///*2g4<aeWadaXegdVZdgggp����������pgg����g�pg��g��Ǟ�gp�gmea<32/*23X/*22V<<aXgpq�����pmp�gaaXVa9/*/*//0<22959322/9<<<95<<V<XW<<352<<<5XV`999227///259<XdXadbWefe<[dggfp����������pgg����g�pg��g��Ǟ�gp�gmea<32/*23X/*22V<<aXgpq�����pmp�gaaXVa9/*/*//�XaefgbdXaed[ep���p���ggeaX<959WX<VXda�qaagmeddV2959Waea����dmp�m<X<<XaXegp�����pm^V98////3<XaXXdX<eaXWagX<<XWV<<233252/+/+53<3<X<93//392/3295<WX<[XaegfbdXaed[ep���h���ggeaX<959WX<VXda�qaagmeddV2959Waea����dmp�m<X<<XaXegp�����pm^V98////3<XaXXdX<eaX�X<R<X<<XXaXedXa<<5<523WV<Xp���dXaeppegpg�������Ț�Ș�ǘ���qmdmp������hdedW93mm�pmwmdmddaedgemdaaaefepefedd[eaXaaepdaadaXdaW5W5aXaaVdaXWa[dXgdedXX<5XWVWW<<X<<XXaXedXa<5<<523WV<Xp���dXaeppegpg�������Ț�Ș�ǘ���qmdmp������hdedW93mm�pmwmdmddaedgemdaaaefepefe[253                                                                                                                                                                                                                    9aaa[92
[523
93<<9V�Xdd 


























a�dmdmef�aXa/802/9937979//707/906/70=:9<^?999=<=3679299////7//////062/399078096/077/906/70=:9<^?999=<=3679299<g��mepp�h�[b[0<<XXdXg��q����gp��ppbaa93/3<99V`baa<^pa<9^^V^^ak^bmampqakbka^Xaepmpqpt�wqm��ɲp�eVaeapemdkaVV99899^a<^b^9^<997806979aX^aXaVa9<9339VWVXWV<XWVXWVWX595<XW<XXdXg�������gp��qpaaX<3/0<<9:`aaX^^ed99^a:^^ak^bmampqakbka^Xaepmpqpt�wqm��ɲp�eVaeap��ϲmaaV^<�geg<eggp�ggem[aX^<aVa9<<aaaXemdmdappmaaaapq���pm�wwemvpemdkaaa^dw���v�welbaa99mpema^9<^a06<X^<^989?V7279939<909?V`aaaaV9<8729^`V<V<<<VWaXXa[dX[[ded\mfe[aeggpg�gmegaX`^<aVa9<<aaa^empeaepmelaXap����mp�wwemvpemdkaaa^dw���v�welbaa99mpema^9<^a08a��p^<99<^
�aXa7[eaaaak<X?<XeadpbWbadaX^Xepdmaeedp������eoppwpqw��pw�wppme9aae=V9bdqplampbalaa^a^ama^XWV89<V<V`<^^<<9<V?<=Xaa9V?<V99<99<9<VadelgepeedgpededdaXadXXaeaaedaabadV<a<XeadpbWbaeaXXaedplaedep������mlgw�pqw���w�wppme9aae=V9bdqplampbalaa^a^ama^Xgpgm<<V?X<�XeX
/3<VaXepaaXXaaWeg`edXep�������pp�����pepdme����pgpp�meammqvpbpaapmdamwmmmdmpmwp^aV^XaWV`Vd�pejaV9999<999V<<VWV<<999<399a?^a^^<^<^V?Vjeeabd�emeda\a<<<93<V<XaemdaXXaaWee`efXdp�������mp�����pepele��p�pm�q�mdanmpwpbpaapmdamwmmmdmpmwp^aV^XaWXdp��gmaa^9g<V<^gppepaaXdbdagmpgpp����em�����mm����w������pmdaaaapaamg�mhmgmaaaamvqjakqma^V7^aXe?abdeaaXaeabX^a^<V9^Vaa929973?V?V9^a<<^aaba?aVaaXaaaaaaaaaXX<<<V<VdeggppgpgaaaaeXdeppgp�����epq���ppm����w������qmdaaadeaampqppemgaaaamvqjakqma^V7^aXe?abdeap�ȟadVaaV�aaV 9VWaaaemp��������mmedabdbdedadXagpdeedmgmdmep�Ĳ�����mdpe��mleala^aabja^X?XaadmdaVW^aemppmg�pejelpe^W^`X^aXaaVajX^<a^a<X?aVaXaVWVWV<X^9V?V`aV<eaa^VaaabaX^aaemh��������mmedabdbddedaaXpgemfblgpaemp�������ppepd��elmala^aabja^X?XaadmdaVW^amp���ɘpmblm�^^a7amgmbmlemeaabV^ade`ed�egpd[ep��pep����v�����q����w���e��ppq��qv����wppv���m<aaaaajmmmVaV`aa^a^VV^WXdaeaa^daka<addeeaaX^W9<X<<</<Va^aemoeaaV^<^V?aabaaXampedmmmemaaX^Vaedade�gmgddep��qdp����p������������ğe��ppp��qv���Ϟppv���m<aaaaajmmeam���aa^^V<�^aa7aaa^da^^Xdaaepmempgpppg��p���p����p�g�dj���������Ęmp���ɘpppw�mqppmpqmgbl��kmw�pb`aa=mpqvdaaele?bdeja9<?q�a9aaVaaaX^<aaamWV99W9aV^W^daV<aaXX?aaaampabjaaXab?^Xdaakgpmdppgppp��p���p����p�ppdb����������wpe���ɘpqpq�mqppmpqmgel��kmw�pb`aa^����aaadme�mpm/^agagaapgpeppgp�p�p���peegp��eaadepp���������������eadXaepmp�qppmpelme^ambj^bdmXdeampgmvq�q�meedeaaXVaaVa�la_?a<^<9<Vadada^<aV<^^al^emjaaXdlebmpmmma<9aaedmadeppegppp�p�p���peegp��edaaepp������w��������eadXaepep�pppmgmdmka^mba^bdma[eampp���ژwpede�amm^gpgpgmgmpepdpggpegfp�gggg����p��qmw�q�qepp�ϟ����mdp���ȟ���pmdadmdbl������p���qp��meepaXaVaaa[ea[pdeama^ej^a9aV<?aaa^X^X=VadVaX^Xa:`abWaemeldammdmeepgppgpepepgmepggpdggg�pgfg����p��qm�q��qepm�͟����mdp���ȟ���ppbadmdam����p������p��meg��Ș?Xabdd�edV0Waa[aa\dadXX<V<adgpgpgpd�ȟ��������pp�dp��q�p�������p����Ȳ����pedg�pm�gpmqe�p�pgeddddXaXaammbmpaWV?9///6999<aaab^X^<XaaaXX<X<V<V?d^V?V<^d?V^emaXaX<aXaXadYad[adaW<VWaed�pgpeppȟ��������pp�mf��w�p�������g����Ȳ����pdeg�ppqppmpe�q�pgededdg�ǲamkdmp�a^<<aglXaaaXp�����p��ǲ����������Ț�������e��ȟ��������̲Țǘ�����p����������e�pgepdlpbaeda^aabaa?a^a^a^<:9aXjejeaVXaadaaaVdbdXdaXeaaaa^Vaa?XaV<aX?a<Va<VdeoeaaaXap����p����ȟ���������Ȳ������pg��Ȳ������Ͳ��Ț�������p����������pqppepdlqaaedp���aa^^a^�9a<0`\mgpppegpeggep�qpppq�q���q�p��������Ț��ȟȚ����ȟ��ȟ���Ჟ�pamdppppqpplemgpppmmpppm�eempgba?^aa<<ad<5aVaXlaX^XaX^dXabd[X^W:`VaVa<aX?Xpd^<aV<^<<9<VWaeglg�pegpmgfge�qpppq�q���pq�q�������ǚ�ȟȟ���ǚȟ��ȟ���Ο��pablppgp�pglegpeppmmppmp����qmda^?pV<V<adpepgpfgdaagmdeedpepgepp�pq���������qpem�pamddeX<<X?<^ea�����ʟ����q�ppp�pmdvpeppeapedae�����pp�pbaWdX[X<XaVdaX?X<aa<9209</////2/9<9V?V`aXXV<V^<XdaeledpepgpeoeXdepdmedmepgdpp�p�p��������qpem�pdmdaga3<a<<^ea�����ʟ�����ppppq�mlppmppeapg���䘞��pq�bda0Wa[Xa[XdeWXagdaedgp�ppedgmppV^<<3<X92/7293//<aV`q����Ȳ�ɟ���Țmkaapv�����ɟ����e���q�papgmae�eaeaaWV<V`V<a<aV`39?9<aV2083X<23/29593<<<a<aadadedX<XdXWdXd[eWXagdaedg�g�mgdgmppV?<<3<X92/08<3/<aV?����ɲ��ɟ���Țvbabpv�����ɟ����m���q�����mXm�mdd56<
/5<mdgpfgp�gd[defeogp��gddXWXaW<XddXXW<<V���������g�����Ȳ�Ȟ��������ʟ�qg����qpgppkbablemfpeaWaaadX<abaelX939895<<5V<992*/2/3WX<Q<W<93a32<95<3929<X<<5<Xjepgfgp�gd[edefepp��p[eWXaXWVWddXXW<<V���������q�p���Ȳ�ɘ��������ϟ�q���q�ppqppbbam����veaWaapV<9
02<<5<<Xa\dXVagXaea<<X29<WV[ddaeeaepp��p�p������������w�Ę���������p����ȗppdddpaXeW^a9a<aae<9V`VaX^aXWaaaaXaedfaXWX<<aed[aeddXX<<32/3//3/39<<V<93<5VX83W9<WVa\dXVagXaea<<X29<WVd[daeeaepp��p�p��������p�����Ğ��������qp�����pppdedpXadX^`<mp��e<9V?Xd<5<
 
//29/36<339239<5<X0VWmgmedeab`<9Wbdagqvep�ɘ������������pvp������gde[d�f�WXXX<9322<<aa^V?aaXaV`aX^<V<X<<X<<daXW<Xa<<5<<<<939aaVX9<V83WV<83832<95932632/292/3<9392395<<X2/<Xmgmedmaaa<9aaeagqpm��ɘ������������vqv������gdedd�f�WXXW<93429Xapp�qaaXaW^�<aX9W^W^bdapedaXV<<aaaW9<:608<<2aaba<V`�pqɲ�ȟ����ppqgmpdXdp����p����defeggfpgXaXWa<<<V?X`Va<eddaa9<<V472<9VW<<<9V<V<95<V9<3/3<</5922<593`Wa[X<W5<dXedaadaVaVaeaped[aV<<aaX?5<=063<<2aaab<<X�pwȲ�Ȟ�����mpempfadg���������deoeggfpg[aWVXX9<<?ag���aedaa<�WaX /9aadaaXaeaV?e<<70/969<99Vma9ae�e^X9aV9a323/279<83aaa�e?Va`X^<Vag���pgogaXX�gafq�pep�Ǟ�dgdep�daemdemdea<d<3///3<<XXaV<3859<<<32W5<59<5<VW9V[bgWaX`<<XV<aadaaaada:VdV<606979<99Vma9ae�mVW9b<9a9323/98999Xadpm<Vaa?XV<am���ggfgaXX�gagp�pep�ȟ���fp�d^ed95<
<93<93<9<a9<aXela^^a`eaappbepmmpV`pa<38VWmd^daXaX<X9/7////V<W^pq��������gddegdaga`eeaadded[edepggagpaXdae[deaVVW93232<952<9X<<XV9<V59W<9V29293<<<3389<<3993<9VW9?aXema?^a<eaappYlqemp<^pa<92VWeaaadXaWVX9/7////V<<am���������gddefeaoXadmXp�̲d\defp�<<X /3//8<99<789/a^a<7////2///<<Xp�p�q�pge</9<339<paaaep��pWXaXaV<<:fepdeedg�����e�qXaXaaa<abdaeddaXaeaapddXaXW<W38<<V<<?X<<<<3<=V<V<<3<3<<<Xd^V<3726//8<9<9789/aa^<9////2///<WXp�p�q�pgb<29<338Vpaaadp��paWXaX<V9<pdgemdeg�����p��̘aaaVaX�<92
295aXppw�qmpmpmba<bppagdaV89<<92Vadmap�ndX99Xepgp���Ȳ��ppeleapd�q�p�medpedaaXaeddeeddXdaae�mdaVaXaXXgXdXXW<<X<X<<3W<VXX<ae^X?:WaXa9W^XaX895<`<32//*2<33<Xappw�wpmmpmba<empapd^V859<92Vddmap�mbX<9^dpgp���Ț��ppepdapd��p�ppdbpgaaaXaedaedgdg�Țd�mda^�WaX 7<<3Waa<//39<<9<**/9<39<<V59/3X^W9V`V<X`ea��gpmV<XeWmdaaemXaeep��pXoXdd[dedge`XdXepX?X^VWVX<<aVaaaXXX<W<3<9<32923899<<<<<<WXX<<<<<<XXXdXaaada<<3aXa<//2<<<3<///9<38<V3<903W^X9<XaV<aedq�eqlX9Xe<mgaaemWaeep��pXp[ad[dgdeg��̚epX^W^e<5<Va2<V9WaV8202<a<99<3//3///2939<99V?X9V?3/////8^999<935////79aam���eaVW92<WV<WX[XaaadV<<aV?Xa<a<9aX^V<?V<Vaa`VaVaXd<<Xa<aXXVa<95V;V59<Xaepe8<<5?b<3/82Xa<99<0*/2///2939<9<<^X9<?9/////8^99899350//99bam���eaX<95<d��gW[Xaaad<95/3;<V9aV^<V?^bW022<525V<2938/929?97m63/63/9<<^99<a<V?<937223//V<7/7///9/7aXde`W5345WVdg<<<eaaWbXa`aXbpeaaXjddXdba<<aaWV<XX<^^9</99//<9<3<<9582///*3<9<V^<^V<=aaV223<423X<3729/<39?97k80/2733<?V99<aVV?99372///20/<V7/7//0//7aade`Q<Qf��Xag<<<d39< 29<dpe<9?:8//02///95`XdaVp��b<2/<9<aeedggdbdba3<8/0/2/6<<[W\f�fggdggaVdpaXaW<<^X<a^<aVaV<<aedaXeddeddaVaa<^Xa<<79<9293<W<<3X<<ape?9<^2/062///3;Xad<amȲaV2/<<<aeedggddbda3<7//2//<WXWg����g[ggaV�e��<eppq�q�lgmaXa?V3a<aaVWaeaX9//22<d^dmp�a99039Xjaeddpp�wmjae^3?Vaa9<aV<e��ZXfXW<3/3<5<<^<<aa0`a9<WVded`aXX`XVadaa^aX?XaXeldbepgdedpg��legdmgo�pq��mpdaaa<V9X<aaVXaeXa</22<d^dmp�a99765^eamddppw�kmada0V^aX9^a<Ve��X����<3295<�dmW
/2934<agmgpdmaepeleW<3383Wbdelpmbdpedba<agpa9m�\</9a^gp�pppe�wwm9<V^9d=999779//9<:amXaaX9<<9//*/23<95<5<3/95<adeaaa^Xabdaaeaaaaba9apeX<XdmW3923</383<5aglgpelbdpmeeW<9383<edelpmeepbdbaWaepa9p�YW/9aalp�pppe�wwm99X^9e=9997736/2em��Xaa<<<
[<<V <dddede�mdXe�baeoVaaVmgaaV?^<^aV99<V/9<3`a9<V//9VWblemaV<//9<9V^9/7Vaaam?^^^<<bda^9^a^V`X:<8WW32929<<<53//0/099<9//9//0*20<<X?XXafdedded�eead�eameW^a^epXa<^^<^aV99<</995`a99V//9V?eejeb^</
/9<9<^9/7<^akm<amw�mdaa^9^g<ae9Ve<<aea<99939<<79<<72//^^ea^a?aem�a��p<<pX^<<<3X?aV0293aep�q�wk���538V/6/606//9<97>?^9<<ab���p��eX<99<?//////3<392/2/25<2<09;3659<aga^beaadV<aea<99999V<89<<9///^^ma?aVadm�a��p<<pX^<<<5V<aX603;aep�vwqkp��539W/6//76/7XW7<:6^^W92/ /<99^<<aV<aa^aVaX<Vle`^X9=V<93<<29<98aqgmdmpp��vqpggedaeaqa93?0<9<X?dedaaam`^ml:8<9V<V96/9//990/3//////3<<2809V<<9a^<9<<3/<2///0<99^<<aV<aa^XVaX<Vle`aV<9V9<9<<09<98ahpmdpmp���qpeggdbdbpb83^2<9<^Waedaaama^ml><9<<<Va^de/p3`a
/79:99/39<V9<//23W<a�q��pbpm�p���qpmapa3/9a923<3<9V2/<aa0/7//92<^<528Xeaemla996ma^<?9^<V<<a<XW/8*02/3/*5VWV^a9<0///83//3<<89V<8Xa8<ab<99?90/39<^59223W9d��p�pbpm�p���ppmapa3/9a323<939<329aa0/7//839aV429Weaemla987maV?<9^Xde��<XW/
pV<d9699?3/22/<5Xd<WX<VX`Xmp^3779?0/3W^aebleaaX<<aa39dpaVWd^292<aV`^jm^<0*2/293aaaa9Vd9/ab<990*2/9<9Va<<^93<a9<aaeaaV99/>9<9/22/<5Xd<WX<VWaXep^970=V6/5V`baemea?aV<aX<9dpaVWd^283<^W^ajkaV6//XW0283aaa9^X9dVabdaeleaX<a:<bp�^Xmepd<<dagpdVWV8<993<<0///02/2<W<09dpg<<eaa<9<///792a^699aafdV<X97/^93//<VaWjX72993<<93<VW9/9aV?:?9//299V69<a^XXedea<bdaeoaaX<a:<bp�^Xpkpe<<ddepdVWV99939<<3////9/25W<09dpg<Weaa<9<///639a?099aadgep�m//ga939V<729<<<<<a<VdaW<<5283^b<593295abm�qpmgeav�m�pge[Y</<a^^99ampp^ama^��ea9^XaX9aaV?0/<932499<?<<7<<<9a?79996/3<729a9`398<7<93<2/9<^5<a9326<X9<V=327<^<5^WV<e`X<<<238VaV58323<abd��pepd^w�m�pgdeXV/<a^^99ampp^am^?��ma<^XaXa��q?7/<9d<da7<aeda^X^^XmeW95Vae`Xp�b<apqdeopedaemq����m?ea^<8<X99aW98<9baa/0/`bdeȞ�vemmeamkaeaam^///*///9/<639ed^aV<^99VaX^aX?<380/62/93;9//8V89<9<3<daaaemjX^glaX^W^aemW95VadX`p�a<apqedpppaaemq����m?eaa93WV<9a<<9<9baa/0/`bdeȞ�vempbammVmaam^<<\<//082
g9WV ^<<V<a9?V8999<9aaV<aVa<aaa^<^dXapa9aa938<VaepeXae�madm^^<9^^/9V989/28997299<9^5/2/*/*////83/9aa`V?<?<<W9//9<<3X<X<99X<ba<mp<<<V`9^<7999<V?aa<aVX?Xaa^<^daaga9aa938<VXmpeXalqgaama^<9^^/9<998/39890/<9<VmdX52/*/p09<7<aaagpedmppmeplV?:?a���qalbde^`VaVVWag�edepdmW^83<X?X?<9699/7//6<7daaa98<<3/5269<9/9V6/</2/<53293/29999080/38VaV<9<93^29?<39<aa<aX^aaagpedm�pelpe^9^<^�p��abdmaX^aVa<XWpgedgpdm<a38<V`V`999906/06<7daaa98<V2/3V;/*;3X629
/9<X<<X<<V<V<X99<d9X?<V<Va^lakajpe�apd^dX<Va<Xleaap�q��mak^p^9a</Vaa^=^nwpk��</aX<3//9/3?VaVaa9d^3<V83V9//9989<<999aj^e`<9W^<XW3929^380/2/99<3V<<VWV<X<<V<<VX99<d9X<<V<V^ajakajgmpemdada9VX<admaap��p�mbjkmX8a<Vab?=^mwqk��</aX<a<d<//8V?p<9</<<<VXW^XX<<<^<V^<9aamX?999V9^<99X<9<9aejepp�ep��w�t^mk?>jjaV<9<?aggaa:9^ta<20/9<V7<V<<:83959//32//69X?Xld:9<9<9^d:7=<996<9?V893///3<<V9<`VW<X<<<XVWaVW<<<^<V?V9`bl^<<99<^<<99X<9<9amagmp�ep��w�m^mk?=kaa<9<<^`gpeV?9^tb<20/9<:9<eg�e9595</g<X9 0<<9399<9^<?aX9<^9<999953<58<338<<<apvmlmeppvڟ�w�ğ�va:mele<X<9<?a?m^jmb^W:<aVabaaaXaV`bdVWV<a<ae`X`<3<<2</2/9259<2XaWeme?Va^W<dm<5<VaW<a<a<<9WV<959<V?V9839<9a:?aX9<^9<9995959<3<932<?Vavpmlmmpp��°��Ğ��^^bledV`V8<^`^m?bmkVW9VaVabaaaXaae��ga<<^<Xd5* 2V?^999Vaa3<<<9X<9<aXW9<XX<^W^XaWa^a<epb?dbaa9<V59Vja^dmjm9a^lpdpmmeW9<VaeaedaV?mX<<adadXaaaagXX<aVagaaa�gea9*/2///99*32/3;3<<95<9<WX3259*23<38V<a999^bW9<<<:W<9VaXW9<XX<<X?aXa`^W^dqa<eaaa9<V59aaa^lmam^^adpdmpmeW99<dbaedaV?mWV<ad����aYagaW[Wad/9V<X?V2//9<99<<5/<9WVV`X^WX<<pedbaaXda<<:590<a`V^aamaVaX739X;989292<9/Vd<3239//9a^b<<90938039///23<<<<V<9adaWXaX<<aV2V<99<<952/2/552WdXXa[XW<V?Va<3//8599<<</<9WV<aX?XX<<pedaaaXea<V9<90<a^W^VjeaVaa363a98989229<VdV2229//9bd��e963930g<9<
 
2^<<<pddpdep`[aaa[W<adaaXXWXWX`ed<paaed^da<9a�mam<daWXa<<5<W<<<a<2damV?ab`?apaemaa980998=//45WWe[g[W<V39<7p^*//3//2<<<3;VWV<<<X<929<<59<9594/3<<<<pdapelpXdaWadX<`daaXWWXaWXmdVoaaedVda<9a�mam`aX`Xa<<5<WW<<X<;aXp^ValV?apaemaa9Xoa99=/pedd7aadaV`a\a<^a[aj[^<ddX`XV[dpppeda`elm�vdedpejaaaepmdbja<WWdlm��������ɲ�ğ�mpqppabdgp����mp�qmaWaW<a\aYaWa<<5<<<^9<92323<W3W9<<593///3<5<W/<<VdeddkabaladaVaXdd<VadaadV<ddXaX<[epgpldXadmd�wdlepdakaadpmeabj;WWddm��������ɲ����pm�ppabdg������ϞveaXa�aXm99Xad\d��[pej�^<a?�e?X?agp�ĞpXdm�mapmeaela^<maam�ğk�������Ğn���w�qqpqpm��eldg�gpemdgeaaka^?aba^VaV6/22<39332<325<W5X2232<<92V<<V<<<V`V`VWaXaWma^<9aVWad\d��\paep`Va?�e?X?agp�ĞpXdm�mjpmeaeda^^djam�ğj�������Ğn�ɲw�qqpqpm��dmdp�pgeelg��Ȳb?^aaa�dX?9��ga<aX^aaWb<Xde�pmppelbjmm<?b��vpfeo���ȟpdm?aw�ɲ�ʝ�ȟppm�qeeaaXamdkamVaaw�kjb�^^ak^9a9^pV?<VX292WdV<X[adeXada^WXaX<<<Q9VaX<bdaaaV?9V<99?aaeaVlmaae��pa<aX^aXaaVWagppmppmdkjnd^?b��vpfeo���ȟpdm?aq�Ȟ�ɞ�ȟppm�qeeaaVdmjbjmVaaw�mak�j^amme�l^pV?9X�aXa9VX9^<9<29a9V`X<W9Xag�mglamW^pp���p�peXX9a�p�p��pbmm��w�pmgeeemmv3q�mmpmt�we����mX:m?^<<5gWV<aX[a<aV<V9?a<9^a`>aa^X?Xa^<XV`<3252<599V9V9<9<^WVaX`^eaXXaXX9V<9<99X9W^WX<<Xag�eplae`^pp���p�p\aX9a�p�p��pbmm��v�ppgbeempv3q�mmpmp�we����mX:m=a:Zp�VWXXaX�a<< 
/?<<Wa<X<Va`Xaegdmpempɘw�wp��pabmdb`ppq�mpq��k��qam^`b�mg���p��V�eppe?bpaa[aaaa8/X?9<<X<^<^a9a76Wa9<9^aba9<9////:</93<VWX4<[d\aXadagaaX`a^WV<X`<089<<<Wa<X<<jX?degdmpempɘw�wp��gaamejappp�mpq��k��mke?ae�pe���p��X�opge?kpaaXaaaa8/a<9Vd���?V^?a7�9<59W<X<5<<adam�pfpp���maev�pmX<eaqmppmɝevmb^<X^a^����ڞ�����ggedaedXjqp�papaXmjb?aa?<^V<Va?:?ke^a?93<V<993<93<<39^W^V<980////39<29V<aaV3<<X893V?<3<<<Xa[?XW<95<adam�pgpp��pmae�qppV<eawevpmɗepmk<VX?b?����ڞ�����egedaedXbvp�gjmaXmjb?aa?<^<<e��m>lb^a^
�[ad<df\dgdXdgeaemaeeepXX^gemmam�mbpmpmp�Xada�gdbadVea<eWggX<WXaadbpea`X`X^<addakdĞpmde��<Xaa<//<5<9<<2<5Vdped9`V92799dV<dba<9<22/*/2/5XWd[aaeddXd[egfegdg[gdXdgpXbpaaegmXXaeemmapwpbpmppe�a^ddppdeaaVea<eWpgX5XX`ademga?XaX?V`dddblĞpmde��Xl��e//<
�9X<
23Wa<WXapdpgddXX<edaaapeledaaWmaapp�ejgm�aVmdea<aaaXba`<<V`^apaVa��q��w�w�v��mqlbX?<<X9?aa9<;<<WaVmgWV<5/3<9/389<</9<9W<53223<Q5X9VX<<<V<X<3<3Wa2X`VWaXpdpgddXXXaea`apeleaaaWej^pp�ejgm�aVmdea<aaaXdaX<<?Xabma`^�����w��q���pql[^X?VW<k��o<<<<Wa�WVWaqde<<a<epaVa[aX`dedade?X^Xaap��mabpabd<abaa<<WdaXaWpg���m��m�da9XagXaV9Va^<baaeaaaVavkaalbfp�p<4385<<X�dge��mde�gpgpXa<aVX<83/389<<<922223;3<X<XWaadm��ed<<a<epaVaXdX`ddeade?XaXaap��ejemade9aaaa<<WeaX`Xpgp�qp��m�d^<XXgXaV:<a^<b^aeaaaVamtm�Ϛep�p<5�ade<X<<W\Xa[aaaVlddedWVamd�mdpgabdabamdep[pWVWQXgp�a5/2392/3W^3<<V<XXddammpkm?mdb��eppaV<a?9<<33<9?V<3<23299VaVW^999?<V939<<<X<abaabaaaaV<W94<3adbde`[<3<a<5WeXXdaaa^ddagd<Vdma�mdpgaejabamdegdgWVWRWg�gd5//3</32XV2<VW<VXddapmmmm?mde��epmaVWp�pd<<39<<�bdV29<<^WaV<amjdaaaaX��ppmmdXaXVdbaalbp</2/2392/1/23<9/3822a49<�qp�gp�p���Ȟ�pp\WdX^`XX<^qa<<WadaV98<949a<8<<994<Vdba9V<VadaVX<?a?0879/0/95<Xepd[aeXaefea<<V?Xa<<amjdaaXlX��ppmmdXaXVdbaadb�9/2/239*/2/1/3W9/3822a8<3�pq�g�p���Ȳ��pp\WdXa`XVW^���pWXdd99�a<a <adp�eada<VW9<V8dX<<9a3m�mX^aqp<<WXW�ɟ�pmm��f�˚g��m��dapl�qvppw��qmedXaaa<X?X<W^XpXaXpedXaXggpeaXWXaWXWW<aX<<<9//329<32/29293<292<3WXWaepX<<aX<aeap�gadp�aeaaX<V<<V8dXV<9a3m�mX^app<<aWX�͝�wml��f�̚f��m��adpl��pmq��qpeeeWaaa<V`V<X?Xp[aY��̕aXggpgp32V9edX^`ddXdm<mqpbdaablelpaV?aVadpp��p�pkv���pmgphpg��m���p���Ĳ�Ʋp�ppd[dagpljXaddaXXcaaXaX^ba?<?XaaX`^X<a<95^XaW<W<<Ve5<W293///32<V<?V99<93a<93<elgXdgaaVaddXae`mpnde`^dkdmpX^?aVaeog��p�pbw���qepe�gp�vp���m����ğʰp�ppfadXppdjaaddaXXacag���aa^<?Xg455<V`emeppejgp�qpppaeppmdp��pgpqp�pmqp�ekgvpeaXebdaXajepmaddaaXddebdbpp�ddaadbaaaaaepdedmde`eaXaae[[dXa[adXX4939dbd9V95<<3<98^<9^aV95/7<9XV8X<552<5<<aaXmelppeappq�pqmaepplep��pgppp�pmqp�dkpppmaXedeaVaampeaddaaXdedebapp�dddaabada?aepdefm�ȟ�aXaadYQ/2
 <mp93?=pa<X<;/9^</7W?9^�w���p�ȲmedeWXdf[a<^aabd`aamaamlemddpdaaV;aedba�?dalm`Xa`egogaXeddXXagXa[a[XWXV<a3<aa<aaXaa<^<<?99<^^9365<Xdd<2<V<32**/23?a<mpg98^9pa<W<</9^</9<^9`q����p�ʲele[XWfd[a<^a^ea`aamdammmdmdfd^a<?ddbabpaadle`^dXdpgga����XXagXdpabd9<95?a��Ęup�paeppda���ɲ�ɟq�pq����ȟͲ�pp��qaWe5Xdgemlmpmppdlkmmlma<?9<Xaaama`aXW<XdeeWVaX<XWV<<<<<<9<<ag`///9=939<//3//23/9<9<W332+2+/a<<daeadaae<9<Va��Ğqq�maepgla��ɲ��ʞ�qwpȗ��ȟϟǘp��pXadRWdgemlmpeppdlkmpapaV?9<Xaaama`XaWVWde����a<WVWV
d/0 /0V?3///29<Xee�ƚ��p�pb<99^e<Xabm�������e`d[Xddkjm�Ͳ���ɞ�pedamg��dXaXddXaX<X<X<990638<9<amaZde`XaXdVXapa<aa9?deg?<a<<X9/*/2V<9a3/080273/27/09<9V<92/2<<Vdm�Ȱ��p�gaV99Vp<Xakm�������mWedWeamam��ȟ��Ȟ�qdejdp��[aXaddaXa<X<X<eaea72<<9X[2<<

Xa<<XaadeWpb2/38^apwpkmk^mma:9<X^����pmv��v����adedXXW[a?<33<ZppdaXaW?epaa�mg�p�dmdXe�daXW<<5WbaXlXadae`aadbd<<395<Vdp\m�b<V+2<W9292<<////2XaW<WaaeaXmd5/92^avqpkmk^mmb99<Vap�ϟpmv��w����aade[XWa`V<32<[�padXW`<epXa����͗gedae�dX<<Vdd<jg93<X<?WXaX9XlaX`e?3/87/<3<9���������ɘp�ϟ���Ț�������ȟ���p�p�ppppadeededped^`Xa[aeal^VlVa<aaX^9^a^aX^X9^Xae<932022Xp��epaXWV`X�pXdd9em8/3<X<<aXaV5Wea<ad^9/9//<59<q��������ɗp�ϟ���ǚ�������ɟ�����ėp�qpw���\dbd�ee3<d 
7?aVma23///=�kmmbea572392<^8a��a66<�9>89/9207q^^abXepb�������������İ�����wmm�mpmqm�mdedegmdpgmd^lV98<<amaaamo\dbp[gdaXXabdada<<<<<5<3<aa0/83<dXgdV99^`Vkd02///=�kmekea<02992<a2a��a/6?�9>8<33/07m^^Veaepb�������������İ��²ɝmk�vnpmp���Οepedpm�<23/lX9223<lX`aaV//5929<edm��gv��ɲ��wlama/3/3//3`X<9apdb������xm���Ȳl���ȞĲwq�����pqpp�eleemmplepmdeleldeaadad<aW<WV`XaeaX</93<gaX?aeaaV<222/2/<pW9323<lX`aaV//5389Vded��pp������vmam^//9/3//3WX9<^�ae������wn���Ȳl���ȞĲwp�������gp�mde5/2W

2<WX99kmwm�mw�mmXpp09da*/*/<VdeemXbjqmapk20/7^lm���p�mmqmkmVpVaaepmp�����������pqmdppgablbadmpq�q���pp�goXaXd<9aaa<a�a^aa=aa99/+2<<5<4<XWa39kmwm�mw�mmXpp39da/*/9<eedmVblpmbpj3/06^mm����pmmqmkm/5pVaaepmp�������⟘�pqmf/2</2X3/////^a9////2/[X<8<6/^a8V��͞ppmmpa2//*aa7^=989Vmdadbaepep�9dV/2/<VVbaX?592V<993<Vampea<^^<<9?:a99<?a?9?9/2<2/<<<<2/*/8X2*////:j<////22X[<8<6a`7W��ɟmpmmpa3/j^9^=999<meaabaepmpq5aa9V^3///<g/699993aa<*4e`<p`aaema?^937/25<3a/679^�madbd�V</^elpg8k?=7jm=��maeW70*/X9/4<<?996/^6//2//699/99///99<V/893<7<aV?9?<<9/89<<^da9<9VaX5f^Wlaaaepa^<990/25<3a/006^�madbd�?<//?empg6/k?=7jm=��madV90/X9/2d�f^896/^
a7?/ *8am��Ęamka><ap?956069a<9adk99=^qm<3mbɲkvm99//6a<d^a�lVjmajkadaampĝd`<dalppv�e^=^ka^<0a60/7299?ab`<9a^^9609V69V6*8ae����amka><ap?9<6069a<9adk9?9^qlV2mbɲkvm99//6^<l^a�l^p�ɞkadbal�vea6383<a�pmmk^=k��wϟba/6ba<9Wa�