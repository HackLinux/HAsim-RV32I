hanges you have made<br>without closing the Java Control Panel</html> ]<html>Save all entries containing<br>product name, version and<br>location information</html> .<html>Save changes and close the dialog</html> @<html>Search for an installed Java Runtime<br>Environment</html> r<html>Select this option to show Java<br>cup icon in the system tray when<br>Java is running in the browser</html> T<html>Select when you would like <br>to be notified about new Java<br>updates</html> R<html>Show Dialog with Exceptions when<br>errors occur during applet loading<html> '<html>Show the Java Cache Viewer</html>]<html>Specify the amount of compression to use<br>for JAR files stored by Java programs<br>in your temporary files directory<br><p>With "None", your Java programs start up<br>faster, but the amount of disk space<br>required to store them increases.  Higher<br>values lower disk space requirements, while<br>slightly increasing start up times.</html> F<html>Specify the directory where temporary<br>files are stored</html> \<html>Specify the maximum amount of disk space<br>to use for storing temporary files.</html> )<html>Start Java Console maximized</html> )<html>Start Java Console minimized</html> R<html>The Java Cache Viewer cannot<br>be shown before the change is applied</html> P<html>The Java Cache Viewer cannot<br>be shown when the cache is disabled</html> Y<html>Use Sun Java with APPLET tag in<br>Mozilla or Firefox or Netscape browser(s)</html> I<html>Use Sun Java with APPLET tag<br>in Internet Explorer browser</html> 4<html>View and modify advanced proxy settings</html> H<html>View detailed information about<br>the selected certificate</html> ;<html>View information about this version of the JRE</html> <init> 9A mandatory update is available.
Do you want to continue? About About - Java 
About Java About Java Plug-in About Java(TM) About... /Access to persistent storage denied for URL {0} Access to {0} failed ;Accessing keys and certificate in Mozilla user profile: {0} Add Add missing root certificate LAdded SSL certificate in Deployment permanent certificate store as alias {0} 8Added certificate in Deployment denied certificate store HAdded certificate in Deployment permanent certificate store as alias {0} 9Added certificate in Deployment session certificate store ;Added certificate in Root CA certificate store as alias {0} ?Added certificate in SSL Root CA certificate store as alias {0} Added progress listener: {0} @Adding SSL certificate in Deployment permanent certificate store 9Adding certificate in Deployment denied certificate store <Adding certificate in Deployment permanent certificate store :Adding certificate in Deployment session certificate store /Adding certificate in Root CA certificate store 3Adding certificate in SSL Root CA certificate store Address: Advanced Advanced Network Settings Advanced... 5All rights reserved. Use is subject to license terms. Allow JRE Download Allow if association is new +Allow user to accept JNLP security requests FAllow user to grant permissions to content from an untrusted authority 1Allow user to grant permissions to signed content �Although the application has a digital signature, the application's associated file(JNLP) does not have one.  A digital signature ensures that a file is from the vendor and that it has not been altered. Always Auto-Download Always allow Always allow if hinted Always allow this action. /Always allow this applet to access the printer. 6Always allow this application to access the clipboard. 4Always allow this application to access the printer. )Always trust content from this publisher. �An icon will appear in the system tray if an update is available. Move the cursor over the icon to see the status of the update.  IAn optional update is available.
Do you want to update the application? 
 Applet FApplet supports legacy lifecycle model - add applet to lifecycle cache Applet {0} {1} Application Application Error Application Update %Application unavailable while offline Applications Applications and Applets Apply )Apply jardiff for {0} between {1} and {2} MAre you sure you want to completely remove ''{0}'' and all of its components? :Are you sure you want to remove the selected certificates? Ask Me Later Association Warning GAssociation already exists with MIME type {0}.  Do you want to replace? GAssociation already exists with extension {0}.  Do you want to replace? At: Authentication Required Authentication scheme: {0} Automatic Proxy Configuration "Automatic Update Advanced Settings 0Automation: Accept optional package installation Automation: Accept printing $Automation: Ignore hostname mismatch /Automation: Ignore untrusted client certificate /Automation: Ignore untrusted server certificate -Automation: Trust RSA certificate for signing EBad MIME type returned from server when accessing resource: {0} - {1} FBad version in response from server when accessing resource: {0} - {1} Basic 3Bean cannot have both CODE and JAVA_OBJECT defined  Before downloading Before installing 8Blacklist file not found or revocation check is disabled %Blacklist revocation check is enabled 	Browse... Browser Proxy Configuration Browser settings changed. 'Bypass proxy server for local addresses Cache Size: {0} Cache Viewer *Cache entry found [url: {0}, version: {1}] .Cache entry not found [url: {0}, version: {1}] Cache is disabled by user OCache is disabled, cache limit is set to {0}, at least 5 MB should be specified Cache is enabled  Cache is full: deleting file {0} =Cache must be enabled for nativelib or installer-desc support .Cache size is: {0} bytes, cleanup is necessary GCached copy of {0} is out of date
  Cached copy: {1}
  Server copy: {2} Cached file name: {0} Caching classloader: {0} 2Caching is disabled.  You cannot access the cache. 9Caching is disabled.  You cannot access the system cache. Cancel ACannot delete file {0} since it is being used by this application GCannot delete file {0}, may be used by this and/or other application(s) -Cannot download resource.  System is offline. "Cannot find jurisdiction list file FCannot validate SSL certificate.
The application will not be executed. �Caution: "{0}" asserts that this application is safe. You should only run this application if you trust "{1}" to make that assertion. Certificate Details... Certificate Path RCertificate has been verified with Internet Explorer {0} certificates successfully HCertificate has been verified with Mozilla {0} certificates successfully DCertificate has been verified with Root CA certificates successfully HCertificate has been verified with SSL Root CA certificates successfully SCertificate has failed the verification with the Internet Explorer {0} certificates ICertificate has failed the verification with the Mozilla {0} certificates ECertificate has failed the verification with the Root CA certificates ICertificate has failed the verification with the SSL Root CA certificates Certificate to be verified:
{0} Certificate type:  *Certificate validation succeeded using CRL +Certificate validation succeeded using OCSP 9Certificate {0} cannot be used for client authentication. Certificates +Certificates for {0} is read from JAR cache Certificates... 	Change... aChanges to the next-generation Java Plug-in option will be in effect after restart of browser(s). 6Changes will be in effect after restart of browser(s). Check Daily Check Monthly 8Check TSA extension key usage info failed in certificate Check Weekly -Check basic constraints failed in certificate /Check critical extensions failed in certificate -Check digital signature failed in certificate 0Check end user act as a CA failed in certificate 4Check extension key usage info failed in certificate 