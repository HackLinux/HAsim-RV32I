�6(a@��Ԭ��||��A�I����׵<$����ѥњٚ���Þ+H-aB�X���kC�Ᏸ�x�E����m9a�%���Ӭz��R��I�1k��8z�s\?8E(��F��ˁ�ixm�M-���n�Y�g��|H�������eoÉ{^��f]��G���S���h���t�so�T�oƎ��s�((�V\�Sn7���G�R�ɼ��$�<��nͺ�-߶���D�[g�ئ�kB�Ai3��}+D�$B�b1$LfI�.e��y�����&<d�����z��*�`/�8�4�����}Ҥ�d������A��Y֮�����s�mmxO��ۭ�f�X��P86N�NF�L�,�U�C�d�l�[[�׏6eTTT?��~��,,,���yfggޠ��	���� ^�|�RCCC]]]DD�������$''��qqqmmmnnn))��:::���������}�M� �����WW7"�7"BC{�����{��~hKF������J��A˄���+�?��2�\C@��3�$'x����}������!�"\Y�jר�'|m�HȪs+�mX���h���ږ~8g�a��!�={O��-A.���"����j��n�.���[�.����@bB��T֔��La�hQd$�%NT�C8�D�\BsYTy�EW�%jq_�F��v���H�Z��� �9���_������`u�f���d��������~��{d #��ms���7B�Z�5ԇ�A]a��v},���!�xdGu��G_\��AM~�`�9��_�X��	��ߒ��Do�������e��@z��܅���8����]��WFH���*�簙x\5*�;Ɔ[�5��������Ep<Vp�tԨ���QD���(�oi����Ug�����9r& ��B�`=ɍ)��@v�g�4�������������f�f��9Yg����
T����h
"0���#P�X#�֠�N֟���R ��C�C)������j5����1�3��R�,y��^�J}����w��}z"��i%s-���L�Q��J��9oi��6�2�r|z��`��`��F*[/��_���w������ׅG#~ܧq_��������Cba����*��"�! �ۣ��MY
����C�3$A��o�;����B��u�7jr�AjK;a�ь���Շ\�����&����׷��n��i�_5�-���
IP��t������r���{����3Y�_�v�����������_��_�'����߰�>?auT</�b�qٗ6?153BN��TޥI�+#s�[$���9p��=��t�pt���[�O�;��6#���I:�(B_�B��h������,J�*^A���ԇ��R��·&��HR;���Id[4�p����*/�U�;Ο��CW�~�I\K� ֘j9�ȭ:����8\~�y�Bc��I/0����YUGr�O��x4�i�k�>��<��U�E�3�D+�M)A�yf m�ԡ�^�U��!�ޗ-/Nz�;�R%����+�N7�^��p5��-�Lcp��A�s���9��ܱ}VW3{�Gc����>�b2q����\B�ZF�f���H��k�w\���a��4�N���O��􆽵?�$�hO�+'��]5S���yaU�cAZ.מ���>N��	p���@`D}QOjeߧ;gcF9u1-�&B�����l�V�Sp�+��l57�J��־�bf���3��9Ե�]F�ė�etLQw$�u�l��/������}�u�V�]��Ж�&�MX��ʄ���z�I,�
'��t��+I8�3;��D�v��ν�؁�]�/*]Ì�u]�L��<2I��>���Ԕ����i&G�R�Ab���&f���t�8���f����.k�ǷK:�'t#�ǻ�tQ�������x��%Ӎ8��0�dl�5u���~g��OY�4�YOO����n�Iuv�[_#`�Fm�J�0�u�"�o������|�eM��H�������)`Hs��� �@BH� )QQQ ��
���v&��JJJ?�W����"�p�q� &���ddd~8�IKK	YYY #//�i����QPP ��. ������@BH��W�oЬWWG_����GFJ���,,~@��j+�O���^T����@6w�����AK\��U;�%X�>OG�]�0O�4�[F��F�����B��m������.2�N������`�'Ƴ;s�U��aJQ,�bP%ϳ�-��bP��>tgS�ƘKc�W�`�0�	BZ>�F/V9�Q��x��O����e�ԛ��$��!�X&\�̒�C ���F
���������O��=jq���c�L���_}P��{���{K��Vc>�`#G�x0����d����-���Q�ӯN�Gwz761�}�s���+�+�i׃�*m�t����{$�r~����������K\Sz��Y�9�͓�����h��8��d��t�M�K?�VCU	T{��B=�@B��!o�E� so�����1�|`&:0E�2̡����j�s*��^��3�Xi�ZW�.�l��02���)��(���@v+��� �khܷ?iG'�׎��o��	9�I�Wc��i��gh\�t��e�݉>����d�ü$j\|+���`�.�*���%q�M��׿��H �� ��&V���F�<z	�?9�J��>R0�38���8���p�'p�&���o!]�-34)�(xX#�"�3���@��
��|�Κ)s�mMOJ��2R2Ǽw>���fk�5�;���3*���?n��I.@R
�] 'M��>��%mpA=� ���ٳ�5)1%�L( 4MZцl.�5�C31��6ŏWlw�YO������aɳ_���['��Hp�I��a�D�p	���DBQUv��R��}YN~���i�ے���,�bf���Е-�j�E�̹,v+ƺ��>@j�Xu�6�W|��4~�j�^0h���^�y��2�4�C
�}q,]T �ڇu.[P<%F�h�.�*�73*Se(�*]$�[��3���R���C�70ñU��yj2�e!���%b�WW}�<���\aX"��[/3�%[|��� ����Cq�zF�"uB)��*��5ꦕ�^�y	ik��}��	T!��,ӇL�Fh.E�J��eA˞�E|������(����'S��4]+���Äs�p�
B=��3axD8U�S�1I@��9)aV��XYQn���E2ƪ�;���t4��s/�
������;��)�j��5D*��+@�ۙ_���V�1T��c�z� �bxZx����~7�*���F/����?_>�T��˸A�Gd�]��4��d��$�q�@