.c-Y$_��+OPh;*�"e�b�Y"Ez��j|׻*� �\�'�r�U�ݞ��-°�3Ա��X�Y�ʫ:��ʫ+��2�i*:jd���qN���)N:����S/5)r������O���o�n�q��Ҷ�Ŀ���E?���� �$�|5�~֖	5̓���hgDFJ�K"�f��Z�?$��� �f3��F�v�a1"|��}�ڻaZ�:����ޖ��CFx���yj�u���'�>���m�g�/���Ҡk��_�}Kx�=z���o��\@s�����]"��P�O ���C3�\�#V�8�,�"�����{�4���E�����p�g챶����Qz�=�[����,���B��8�����e����n(��pfrg&ٶ�~�0 ���W���W$�r{ž|6ze���:��!?����qB������l��[����NOg��RAt����V'�ț!�ZWr�Z�x~P�Qhh���Z#2�J?������l���z=iM%�Y�Z#�1�����r��N�O��ܵ�N�]�]T�PM���I�ݠzc�6�X)'�>ZV��;9�� *���m����k1~�%�T!�f��Mz�����(��Vp�~P�=<�7�.YM��ˑ���B`��n��
O%KS��J��X�4a��N}��n�%��\�����+���a��5�C�y H�ڥ8d�S�%AH{�3U��@��}�Ene�%�1qS�5��NfΓ�T,�8 �y�>Y�5M#}>+��S%�&4�/>������Z������T�Mg�j�J?������%�Lʆ��UϢ���-l��b���4?O�I�=C+0[~롫`��0�|��B�B�
�ߊ����wfdv:��9�*��H�lښf�8�����e�9?F�}��&u�������i��!��@uw��P0�� �K3 ��`:{�-u�Y�Q�j�`������t�A���މ<^�_B�oW�5=<14>,[P�,��$� R��0���"G��2�x��R��γ�����:��$���@�Q���zMJҕz��ϧ����Nn���1���PU�/���M7Ps7=Ȟ_�t+n�+��](�G�BD�ռ~�?����H��"ٞR�{c"԰�9B+�"�t����B�L�����l??{��L�fK*~%g���Ki�$o��r��o��Re�"Dr��%&J'f��@S���Gz#�N�gC�kQ*0�1�l���y d��<}e�(���t�r�?1b����pW��rM^YP��W�/(��&��+2�%�T�&bZ�Jd1׊��1�C0 �റ�`�8���@�����9�Sc�J(|r=2�T�����ܖm��Bx��S�"��4����╹U�rVPջ�	�6
��kU<�dIm��y�%O�����Ģ�/�͈&�M�}�w�>��[�R$�@��7t�A������3�
6	3��f�8��N��E�K�w6i���t��ꮚ�fg�5��v�Fl~��m�/�z��1~m�,2�!'���[,}�^��u�Y�2>J�>�Ф����h��T~J�W�R�h�mƝ�ǉ�����a�yV���2��|�}�U�fi}d��&]�dns������b.S��;��Aph���O^��$8(�^�W<���󹶺s�F���C��M(vJ|��\Y�y��P��[�{x����Д/P2�SS��������.���1sy4�,��J��X��X�"T�������Fy�C&e#��<���ͩ�u�;U�oE��=!n�A�L}��рN�'��׽MWI�`�(���&�o&��������B�k�N�N�&�+_dh����y_b�X��ll�q��C'��d����8N$���� ��M+Yl�V���	ϩ�������5�wl�h]���[����޶1�/Y�sC���Պ�PF�FS�%�<�-��zO"����s�ZKf$b����ձ@���X_�8���5԰���o�]�����C�������6]h?������"�A���-w�0igǆQ�l�Wq��P����,e�a��/��:��G=���0/x,�,��!��i��>�f�(m���`u� ��J�������M�1��`x�^��X������RH���@6��va�%S�jyP��7�V���#�%����B_>��dK_�d�+�d_��A�Κ��V[3�87�L���[��2�#�(��a�N8�2	L7���!%��4t������I�r�/�>�-��1O��M���y�&zJG�{��KU��o�Gb��%�_h|Vfk5"�a��uhiKJ�m}��*!U�<�*-Æ	5�y���)�
��),
�pʉiA��b������m������jFW��\Rf���f�*�,+���	$�~�EwV��##�hm��S_�b�x�ݛ/4���� ����_���3��ǎ^���7S����&{a�k�ҡ8�2Z%�h'�Ʋ��v���ё�"�!5Q�P���5g�7�����4ڲ�X�/�Ă{��%��U/)���'M�8V�i�"`I�t�(�\
��,*�*S*����%[*��Db�p	���4����p�SėM��?p�}J���m)�(;�x8!G)�Df�ȯ��	.�!05�%6�H�w]�89��v����y�xP-P#�r`1��[s1UO�$��]6{Kyr��e���u��t����N�Ss1�]}����|�3�۾Ss �{T�{�Y��g ߂��+���$�O7�EB�gJ��W��������F^Y��\|S�