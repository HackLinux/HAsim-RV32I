͋��kDߥR ����A^��B����-��m�m�w�p�e�.~?��xSE6��~��tC��m�L��9G5q����].�����G�g~O����5|fޏՊ0Hh�*q�[Ѝp<�)���$N��-I�掔մ��S��f4x�hzc�*,.�W��e��P��b�e��O����ft�#��f�^Ϙ��)[Փ��S0܄������W9�K`1����J��j?bi���ۋ/\bp�C�I����w5�?0F��P\
3��\�ʔ�/'��A�FQ<`й�rW���n�1���m��UT2LxfU�k.	܊`�ŦXZ�08�q�������C��B 3|㦑��"M�����{Z���A=>�����E�]
�ô�Zz�Rt�U���"6ځ!o�Zb�����q ���yH������^��߁���ޒ�/2WHz���y�T�8������Rx8��xޤ��������Ո<�����j�!M)Ck�v���:@���h@% ��t\/ɀ��� ����9��z��?���T}�;�����)�\-�9��)c	w��|��Fȟ�� �e�y,�{s��ɻ7�P1\ D5g�G�]�� `3A�'Z�:ŢU�� �hM���\� #/ҵ����z�
le�6�HƲ`��
���ML��ɥ	3�`����
 �+�Xa,B/�k�U<b61\u�
�b(�՗����3���^SB
X�f�#�[���+}���kI�Ql�ąv�f��I%�vF���ח�~dM�[�f�2k2�;��Y���D��3$!Ub=�$z�2���N@�&��F���}n,&I�#���D5w_G(��i��H����#4�uVu�!Q'v��#d[�� ����C<0c��C�pJ!'�є��]��(����"�c�2����r�I�"�Z1QN71G�v���(��Mjq���"}��	F�/����pu�t9ë���߀�Du���f���>b&X�>���c���}�i�-m�����ӻ3��n�rʘ��?�br���`9��,�N��ʺz]L���ɡ��C�$��(�����H���,�^"��qg�±��ʻX��m��r��/�����oM��;u�x,�w���:�wL��wL�;�O�ӧ��3��c����Ǻ�w�:�6#�7A�w���>踿�~x�=�e�1}��>�wL��;��[��7��w(�;y�_��L��&�o��������}p�P �]Q�����yɟs�	�I��N�5��׼�_��~y����VJ�?�������\�l�O=]f���F�pfi�h����0�C��y��¿����5O�\Da��/V%?@��N��� f�v$�xp  !T��#�g��f�)
�ZJ�eWh�Og�n��t^��9���k?��Gh������.r�ޚ�[������'�sNӓ1�˼wY��:�!x�q(?`a�}�e`EGp�����P��y�~�;���ܫ�`u���B�=h6�wXs˞c�h?|Xp�D^N� �)@"`�IP�1�=� 
�{@X6V��d�e$�|�s�� ���n@6��'�u:L�Ȱ�᫼ ��"�ռ�:Z��f�����&=�T������ret�@%�ἵ*��,�@��>F ���P�g5��>��ź@S�T	�)���u�8o)`�>/�|w:F�ݲ����F���4r�?�U"��3VWD�t1ѽ�0`0^p`��d'/S��L�Q�_�K*Op�K�U �жVU��ts}	2�58V���;��7ty(�D �^��T6^?a��MTy�i���`���k��}�}�&����2���GBO�4�Vg�����-"�N��T��|Z_-:;���e��|�ï�6�:����G�Ɵ޸��Wz$�O����h�����8�NP���.v��9�&��T?#�G���H���NI����@7�]@��H�c��ʃ�}Dш��߼NKU���aO�3ǪX�:N��Jt���$g���W��?�z�.�*�r4�fQz~�LrNr#�ʃ�dȬq�]]5��c��?�ЙE�R�p�a�^�|�S��zv�!z-<B�~�to�K 5m|����dl��C���=	  ��t��6�J�Es+�v4�����|�	f�T'F��Ӏ��]�	��dʯ�Kk��)�[��8=�Z��_���(���!��<���F�N*-6)N��t��q�m�g��"t���
�'�\K����(<A ���=2�I��?�����-�к�������gad�%'4��"�t}��FZ@>!&JS�#g�����n��τ$7�`�D�>P�����w���k	Y�������F�A�BE�;��%��fqy������)!RZ�J%q�Ϊ�3};!
&�:��� '
f��N� �[�!n)�N]#݉э��aZ���� ��=������U��y��n�x����c0��xL^uP((�d����N����s��&;��z��r����(*E��1��P�Bj��E>��y�/d�8�kǭgǀ\ ��B�y_!!�}�A�)qCnQ*D)��vC'��Q�k���|ԡƽ@�6�`�Ou�	�0�(?�cֻ$˗��	J5�l��yޓ�Q��Y��Q��`�z42K�v�Əm������-7�E�'�|T��i	�u��|�dr�h��2��U���IC��B�p7^�x�2̅^��SK��:py"���t*���U7T;z�������է��R�%��TLFdF�
��mc�طMc��o�kE��m(T�ʇ5%,4ʇ�)���~���Pz�����\o�.�!�l����W���M�U
(�e�1@�ѲD/	�*��C_p<��|�g^ {9�Dw�i1U}�=y��0�&����x�?S���L����e9"&���ȯ��Q4ԝ�B,�u���Qɽ������%�{��t���	[?�إQ��.�_s���,�?K��U��,(�Ś�{9��K�ʹ��=C,���&��q�]��?�)�4��]����7�4��%��@2l����"��G�?��V�@%>�ri������������¯\o�Lگ6��iCȟ�����i{j_$�0~D��b�4�Mj�T7�}힦�I��N�6���.HV�5��y#��Q<�.1<k2�&⦕ϸ,��RmRQG�Br;��o01�R�H�������[e�I�WO�f�{w��G����x�<��zX��*��� $�"�3D�א����͏&�;H�e��Q�й���W*)��_�����KJ�)�%[#�KH�+�b3xm�_���^����K`�zY���f��.��HX��<�T���� �h�%D�秈Y�ĄS��R�9	��e�Rި�E-�A�K@� *�,�Q�F��6��0G� �ș�$��	��Xh� �N��Ž DlR��U�4wQ��P��b�S��D��.[�$�4��E<7�jm`'�Kz$uItW����%v�e���A��e����\���~�����	�8t�	��&�׆>�A�g���rVj)�Ȉq76)�Jʜ��%�o�t�(7���&,Ӏ�1ϜY|���t�k�+,���xZ��k���Tha.������'7����:�)kϰHP��j]@�u�a[�"'�LyrN	��[��15s�%��g���M��-9u�T��T��5���[��Lw�����U�Z�M,���s��'���k��^��T8�����n�C�T_n����{���Ľ�^&�R#)��4�ȱ��Ad88�¼#��q6�W������f�>eh�`��g���S�D}7WD�X�cY�
��}T>)�Ofc�}I2P'�2U�F%'c.;Q����O�|@�1�IŻ�t����|9���p�	�ZS�*����|����f�V�YV��؇��=y��¹����a6xk	qlj�LJ�{��Ke�ś8�Y+'ujV&܈��F�?Y6�nZ��R����3�Z�����#�;m�rs��A��8C5�AC��5�zL�(��/$U���56ؘG���}EXG� �V�n��o���N�k�2_B���+�d�b�xV��jH�Z�U�_?Y�<����'}*����OJ�1��!�o�d�^���֐\$�g������qf��^D��`n���C_D� R:���2ԯ=��H����I~��0`���z�E;��u-�)�ɱ��v
;�����M_�$��<-�"�ki��g�&9��(�}Iz�m1-��@�d�5>�5�Hv�HWvb�!N\]�uԆ��F�(~��.e{��V���كA�61Bi��D��g�R�&�kb-e� O2�Q�K1@q�)����Q������ZZ��XH�m��E�1j�:n+1\�+���+�$��ܛ��¸�G�	4#� �FE��V���%��i����c\��zMl�rh�E�-�F�Ao��<�������,��V+�C-h�ʇ���.�o�d��H��aU�p �o"��3�{�ؐ�����'K��A�C�A��:��X���,c�nI~�srp���{��U^.P�hFZVZ�^1�-PN�A�ǣ��8�~z[�>T6����W��֟"Z{��\�܆�I*ݎ�r���Z��/�f�k��Y�]'���řn��-����e��#H�L������$h��4œ?X��If��)��Z'c�q'8�l3� M(�m��%�W;3���f�D������qhcq���+k��}��4����$�oC�L�+��rF���^;i��� 3�}�秮誜5v��G!�|��^�+��9��1{���r| �����E#����������1cE�yú������	��a��Fz�pf�kU�b�7�
U�d���h@�na3��B|�tt�b�r!R-^v@G)�M�˞�1��]fm˥u缡'.#�2����M��ɾ�����̗!2��/��xia�gm��2 &=q>ゾ�l������s��y�mـ>�a�"j�!]Ve�]���1��'��ز#񚀢_���"�x��4��ʀ&����D�s��&����d��R�P�D'��&�|M(,�'Q�Q��i�Xn'ܾ�+�=ǸegT��ҰW�O���ǝ��蟾��䴔m�X}z��)T<�߫�����=�%\�6Q�^�H��{�Nڈ����*�Y��U�6'�]/��1���U8'H5�2�@���qM���J��fV'6�%
�����Y�]꙲<�]�Z��<l����E�}���[:b51j��wn͏��G�[L� +r���o�^���������JwV�{�C�n�5�-�!��ݏ�n��sp��>/X���llyZ8�rR��H��Ϭ�J���C4���u��_���Zi���	@�)Z~�y  ��wsF�i<�'g���"g��a��o��?SP  ��ߜ��oc8�3�&���&WJ+oז����.�iOf���kx^.����+&>A��"�3��ڐ͈R�Լ-���&�/;�u�zI�)�cN��T6����w�?���m��7q��C���e.�A�,L��p5�f,CJ�Ȅ�cI��7��\�!��3tњ:�'�׬Ǌe��stS ���7�^v͇F�"�mp4��/J�٩�4���j>ƃI6Ňx�ͽ�U����!�ԥ��$�I1��&�1B�o�*��RL_`2䓻�
�04T�a�):�����Ů�Wͭi6�������$�P��oHƃ�������GF�C����C�DE�JY+s�}ş���)�T�d#��h�B���>�b�kf�蠬�6
ؐ:�+��B&�4�a�����?|J/;��g<a���2�c��2}�9�"j����gN�a�j�,�<l���q�m--m�%h�f����jy�M�z|A$H���J W�i��s���t�O�r�q�B<ǚ��Q?��Z��	��fe�ZT�|2�=��ڕ�l~�2;�]�8��!�l8t�H�=7�~�]��ط�J�V�꣭B%6�J��V�����L ն.:9`���R 4X�?�|�2�݈=kV�Nh����F{��G�@�= LZ�'�d�gi�^gm���C�(t`��v��%l�Ž���]�%Ԍ�e�&�gչ��ܢ��®Ĵ�������\��Z�$'��9�/TV��N<Y���i1��[��z�����"�xn�E��`�t�K�\$�R��y��|� K�J쾓V樉�P���#	�E���/�����'.�����=;���ǃ��ΥN?�PX:�\��u�']C�<ć�U�n[ǲϯ� W,�Y�dl���a�1��+��Va�d�d��j �t�bڛ5��Mľ<������Jk���ٸ3��������w�ﺇ�97�V�V�-tv�Q_?_B�.�q1d�ьm7�`[SE5�nЉ?ߔm�A`��`/g=R0̧\bH�,SN���[�-ITJ��+�RD�����b��^���!@�r0S�e��˗�L��$���gfo^�û!�x�_b]�|)?3{F��բ�:���m,��I�@7f��KSn���U~`/�5���nd0��f�o\Vh]s1b��x;y(Ӧx5Dr㦍<�q9Q��i�h���P�<�|L���ε6lh��5k;��C��D�3������D�Pǭo*�4Ů��.y^�c:������I 6�	il��f�