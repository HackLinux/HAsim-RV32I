׾z�`���B<b�S��}��!+���lG}Uo��lFU:���m��Mdz¶�i��>&���vB�i2gj���s`����y]�8�|*���.�v��v#R�D|��ى*�ƺTc���v2��3,||��0,�o	|���g|��B{V��i2y~Q2G���n5�ɾSyz���>e~�G��}��$o��lW�Uq��\KW!:���y��6B����i��8c���vR�D|c���|g����yM�8�|.���8Tj��k*z�8*����|&�˞cc���k1��S0z|��0"�ez���g��0;lV��g2V�I,V���z0°�d0|�ʻD��??��~���$U��mU�W���d:W!:���m��56����i��8>ƻ�km�8*�c��͈z���gg>�|.���sj��v1|�Mz���|*�ˮ�|���v1���BE|��0$lq!����g,��0,mX��gv��;����z ��o;|�ʻ>�~-f�����o��pU�f!+���mGf+F���y{ddP]���i��'N���v|�MzT��͋z����>��*���Dj��k.�yP,i���|&�Ʈ�|���v1���Vg|��0)u�)~���X��I!um��i.���B�|��z4�~@|�ʻ8�3f��~��}o��~f�o 3�|�mW}3:���y:Fb]zƻ�i��'.���k�yP,iN��ȍs���U/d>�|*���.>v��c��6&i���|���s����k&���zV|��,"��,Y���V��;\m��g&|���v���z"3O�E|�ʻ8UU�����}���po�}-3���m:}U$+���m<K+ M���i��1.���c��6&iD�͋|���o)~c��8���6`��ʉ"w�iB|��ύ2��zgm���|8�ƾQl���2-��<,����m2��72z��؋6����z���@h4zMS����PG U�����--���$���QF��̀,G��W:���'f�3w���|*��8>��ʉw�iB|Rj�˝z�����CWv��P���sg��ٍBw�|i���ݝB��zi����P�ˌG~���H7��C4���݀@��H1���ݝM��ɝ����g����{����go4"}��/���<?���4���I{��ڝ9~��y����9��W4G��ݍ6��zB��؍1{�|i�gv�ڝ�����蔔��ˋ��׾����m������Ƭ�����ǒ~����{���p���ﰂ�ǭp������������ˊ���~�����b�lE����h���������q���q�����~��˛�����y���~����z�׾����m�m����쾾����ǏWffofofffoffofofofofofoffofofofofffofofoooofofofofoofoofoffofooffo�}����}��}���}�}����}���}���}�������}uooooooooooouooooooooooooou�u������������������}����J��?!!+!








J��ЖЖ��-%
			





	J���������⭭������oWGLaWGWoxooWUWWeoLaWGWWKQa}}oLWoYGKWfWWWWaaWWWaoYaWUKLWWooooWLaYaaGoqoWLoqqoWaLWWWhYWGOLWooaYWQGGWeWOWoffaaWKULWoqaWUWaGGaqqoLGWooaWGWaLWLW�������J��Ж�������������������������������������������������������������������������������������������������������������������������������������������繦������Ж�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������J����J��������������N���Ʀ�������������������������������������������������������������������������������������������������������������������������������������JJ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������Յ������������J��Ж���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������⵵�������oWWfWLIWaWWoWLuLKKWYLGGWWWoaWoWLooWoWKWaWIWWWoaox�q{�oWq��oooq{t����ooqoaWaou��x�qoxoouuooLGWWYWWWGGIaxoaofhaaWWLKWoaWWUUWaWKGGGWoWWoYaoWLo��Ж���Ж��K-++-+$-	$



����������F3


	

		
		
!
w������������������������������������������������������������������������������������������������������������������������������������������������������������������ǭ����������������������������������������������������������������������������������������������������������������������������������������������������������������{:343-33-3?-3+:-3--+3++-3--+?%-+3--:%--?%-4-+?+--:+?+--3--3+---3+?%--?+-?+4X����F+--%3+--3+-+--%+-:%--+-A%4----+---?%?-?--?--?--+------A>Ж�ЖЖ���������������������������������������������������������������������������������������������������������������������������������������������������J��v���������������������������������������������������������������������������������J�������������������������������������������������������������������������Ӗ���K?<F4-4--34-+?---$4--%-4-4-+-------%--?---?%---%??--+-%------A�����:--3:?--4+4-?--?%?-?-?---?%?--?%-+-?+?%?--???----?--?+?%-?A-?-?+L�������������������������������������������������������������������������������������������������������������������������������������������������������������������������ͯ���ު���Ҫ���Ϊ׭�ҚҰ�ڵɬ���������ޯ�Ǽ��������ڰ�����ڢ�����蝻ˍ輽�~�l��l¸����~��E�m͢S�z��yÊ�қǢ��M���~�b��\�y��yҦ��gˈ��yͬ�g�l��~��c��`����M�6��9zB��B�P��,�V�z9\E��c�m��h�Y��5�E�=Qh�4K$?�;�R��8�B��8����B�6|�Y��i��N�B��9�B��5�9��5�5��0�>�g,Q8��i�9��S�G��,S,�5F$-�)a:�;�D��6i>��6�@��2�Bv�S��z��`�E��P�M��7�,��6�-�|6�B�i	mN��6�h��l�h��2y"�0W$,�)uWC�9�gy�6�N��6�9��6�P��Q�Θ��g�l��P�m��,�5��Bl0�z,�M�r�c��'����MԈ��2E �0K(0�-x<=�5�l]�6����6�dɞ6�g��4�����d����P{@��/l;��M�@�z;�d�|.�v��@����S�i��6I�9<$0�-a4U�0u)��6����6�zŞ8}B��4�Θ��d����R�9��B�7��,�B�z0|g��1�z��M����d�z��1~.�0K)/�"[:q�0f��6�s��6��ƞ8�9��d�Νž]�z��P����B�$��5�,�z"@d��B�y�vd����E�]��6�2�5q(4�,f:x�0���6����5�g֞M�|�ֆ�ΛŮMVP��@����M�)��B{,�z'�@��;�s�S�Y��l�y��*�v�5�/4�)�4W�,�*��5�y��0BNΦ;���ȋ�Ε��EE@��S�s��B�7�|5~D�z6�B��E�`��2����H�w��8�d�5�Y4�)a/~�/�2��5�d��)B;ɥM�v��y�ɕ��Mo/��d��D�<�z�7�|0�;��B�vv�/�3��0�z��5l3�2a45�)G5q�,^8��2�z�� l)ў;ƃ��g��Q��Eo7��S����B�4�z �/�sB�R��8�iv�/�r�)�X��0�b�574E�,�/=�)58��5�4�� \/��9����y�Κ��9�7��l�d��2�m�y'�g�n5�c��#�D�vM�~�"|z��9�Q�69�d�,�M=�)50c�2�w��~/��;�w��g��{l�/qd��M�/��2�7�y8�z�iN�X��B�D�|E���1�s��,�`�5V@P�0�/<�)X��0�Qh�gS��0�/��g�Ɋ��)�E��5x4��"�4vy;�4�v0�g��8�Rv�6�|�'�i��"�N�1hdQ�0o-G�,t5��2�g��s9��/q4��]���4�/|�)I@���@|zW��B�k��B�9�i6}��,�����B�2dME�2�=e�,bI��2�P��y,Ĩ"G@��E��li�9W)y�)K��G1v�?��8�D̘5||i7l/��8�����>�6dEH�0�Cx�0iO��2SC��	I(��$G!��S��BV�C~-l�/K���,�)4��D�P��9g;iBQ*��B�v��96�8�Hd�0�4��0���0�*��h$ğ$U~�G��yg�9:l�-G���1�~7,:��8mB��MV6�cPq6��`�D��	H*�8�l|�7�3Y�2}t�,�P��3ǢF��E��CI�7F$I�$Y3���*��B`P��PsP��;~]vTS�z��g�N|�s5�8�VS�5�-C�2fS~�,�+d�:��Y-��Iģ"7�7fM�4F3��q1�zP96��P�R��;�zvvV�l��M�m���5�8�PP�5u-<�2�s��,F7�	W��O3��G��)<�7fI�3<��	l2��b�2��D�i��P�M|�`�c��/Q-���m�ByzP�6fCa�2~`��0K<�	W��<��4��4Y�7f!I�-<��	|*��M�6��M�`��D�5��P�c��)K+��?7�B�gM�1u8z�2���/Gt�	L��7��7��E{�4Q-=�-:z2��]�5��R�9��2�2��N|8��-e9v�s7�B�;M�1�gT�2�0h�/?)��	=��:��S��~lo\}l\hYoYhYQ\SeIYhal{��g��2�>|�Rb8�4e2i��l�BfEE�2�dR�0�"Q�-W)��	4��: ��4��;749==,;,44-"4#4,--,<;S�i�|.yB�R�c��MY9��<7�@q79�2�BT�04	5�-Ku�	=��$W��9�~SWY_\HIA=YLII70079?Yhlqd�R�|,C/�P؍��N�-��"7-�6f<9�1~,c�,:C��w�	Y+��)~��4��YS;�_HLEGaYl@V9979E�MH�m�M�n	 =v�P�|�D�+��$:�9Y@Q�1�4t�,G!y�o9f�	Y$��"f~�4��S��_mhHEOWq��HM;7=S~���S�0�vgB�P�c��H�4|�m9�5q7;�1z���)�4u�U"��	h$�� K$��3��IlV\lVSQIWlmgHE99SQ\m�ld�m��p�m|�n�p��m�\��7��2�B9�2vY}�}-G�3~�	W��{l�)��QHE\lSMSQLabHH@E9QHh\�qSIE@==9=,4,4=AIQE9E={�)�9�98�1�:h�{-C�G�	Y�� LY�$�~QAElmSVQYWWHMEEEEEQYqrqlhVQLU=GIIC=GYShMHEE��"�5q56�2\(<��-<�	4	=�G	��f)l�-��YGSlld\SYWYMEEEEICIYq�qhqyqqaWYhY\QSYwlhlVS��$�2�;8�*G<�$W4F�	4	B�C�p�Y���SIIhdqdlYSYQEEEEICIYYp{aq�2�qahl\bYbHwSVBqd�o$�9�HB�,C!4�,?+F�	4	E�V2�m[o�'��QIES\wlldYSEEQL@IEIWQqxo{{��qqqdqdlhVdb��Sw��!�9~Yd�,�/4�,<G�	4E�t �mKl�7��WIEQ\wldShSHEWSEQIESQouoqy�m\qqllllbSllldSl��!�9xCE�,}~C�#lG�	=I� W�i{z�9��SIQIhqdSSYMQEYIQVhEIQl}a�lwql~�~y~~~~~~y�y~���6�/0�,fCC�*l$<�	En� L�zO��E��SWQYllSQSSS=IQYQlVSSQq{a��������������������~$�5�9E�,KC�*~5=��n�*F	��#o��=ğYYShodIISWSSISYWmllb\h{{���°��ڰ��Ͱ˪��=!�5�mE�,FO�2�B`��$m�'_'z�6�4��<��qYV�lhSIQ\bYSlYtqlldqbqq�Y֞V�z��nŘ��g�`��Xe$�9�/,�)[Y�8����"G0u�"s1��B�|��E~ly�qlSLhh\~yqhqlllS�yph�D�|1�>��>�c��8�D��6q�9S4;�)L)��>����'�~��"�c��B�m��B������{lYYohq��lYwqldh��lo�n�|�D��>�P��>�N