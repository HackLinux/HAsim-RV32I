cate :Start comparing to jurisdiction list with this certificate Starting applet ... Starting application... Starting installer... Status Stopped loading ... Stopping applet ... Subject Success - Browser Success - Java Plug-in System System Applications System Cache Size: {0} System Configuration System Resources ISystem is offline and the application does not specify <offline-allowed/> Temporary Files Location Temporary Files Settings The CRL support is disabled The CRL support is enabled �The Java Update mechanism ensures you have the most updated version of the Java platform.  The options below let you control how updates are obtained and applied. The OCSP support is disabled The OCSP support is enabled RThe applet has requested access to the printer.  Do you want to allow this action? RThe applet requires a newer version of optional package.  Do you want to continue? OThe applet requires installation of optional package.  Do you want to continue? LThe application can be integrated into the desktop. Do you want to continue? kThe application can not be run off-line, since not all of the needed resources have been downloaded locally The application failed to run. �The application has requested a version of the JRE (version {0}) that currently is not locally installed. Java Web Start is unable to automatically download and install the requested version. This JRE must be installed manually. �The application has requested a version of the JRE (version {0}) that currently is not locally installed. Java Web Start was not allowed to automatically download and install the requested version. This JRE must be installed manually. WThe application has requested access to the printer.  Do you want to allow this action? kThe application has requested permission to accept connections from {0}.  Do you want to allow this action? lThe application has requested permission to establish connections to {0}.  Do you want to allow this action? fThe application has requested read access to a file on the machine.  Do you want to allow this action? \The application has requested read-only clipboard access.  Do you want to allow this action? gThe application has requested read-write access to the listed files.  Do you want to allow this action? DThe application has requested to go online. Do you want to continue? gThe application has requested write access to a file on the machine.  Do you want to allow this action? ]The application has requested write-only clipboard access.  Do you want to allow this action? �The application is being downloaded from a site other than the one specified in the security certificate.
     Downloading from "{0}" 
     Expecting "{1}"  &The application is not allowed to run. WThe application needs to download an earlier version of Java.  Do you want to continue? �The application requires a JRE that is not installed on the system (version {0}). 
Do you want this JRE to be downloaded and installed? �The application requires a version of the JRE that is not installed on this computer. Java Web Start was unable to download and install the required version. This JRE must be installed manually.

 NThe application requires an earlier version of Java.  Do you want to continue? =The application will add a shortcut to the applications menu. 3The application will add a shortcut to the desktop. 6The application will add a shortcut to the start menu. LThe application will add shortcuts to the desktop and the applications menu. EThe application will add shortcuts to the desktop and the start menu. XThe application will be associated with MIME type "{0}", and with file extensions "{1}". aThe application would like to become the default for certain file types. Do you want to continue? HThe application would like to create shortcuts. Do you want to continue? \The application's digital signature cannot be verified.  Do you want to run the application? VThe application's digital signature has an error.  Do you want to run the application? [The application's digital signature has been verified.  Do you want to run the application? )The association is currently used by {0}. 7The certificate cannot be verified by a trusted source. AThe certificate has been expired, need to check timestamping info 7The certificate has been validated by a trusted source. AThe certificate has expired, and it timestamped in invalid period ?The certificate has expired, and it timestamped in valid period 1The certificate has expired, but TSA is not valid The certificate has expired. GThe certificate hasn't been expired, no need to check timestamping info !The certificate is not yet valid. ;The certificate was issued by a source that is not trusted. ?The certificate was issued by a trusted source but has expired. DThe certificate was issued by a trusted source but is not yet valid. /The certificate was issued by a trusted source. %The certificate will not be exported. %The certificate will not be imported. 9The current user does not have write access to the cache. @The current user does not have write access to the system cache. sThe digital signature cannot be verified by a trusted source.  Only run if you trust the origin of the application. =The digital signature has been validated by a trusted source. "The digital signature has expired. 'The digital signature is not yet valid. OThe digital signature was generated with a trusted certificate but has expired. TThe digital signature was generated with a trusted certificate but is not yet valid. ?The digital signature was generated with a trusted certificate. BThe digital signature was generated with an untrusted certificate. >The digital signature was valid at the time of signing on {0}. AThe field {0} has an invalid value in the signed launch file: {1} 'The field {0} has an invalid value: {1} 7The following JREs were found, click Finish to add them AThe following required field is missing from the launch file: {0} HThe following required field is missing from the signed launch file: {0} 5The jar file is on a blacklist and will not be loaded !The jar file isn't on a blacklist @The jar file isn't signed so the blacklist check will be skipped  The main() method must be static nThe maximum size of allotted storage is {1} bytes.  The application has requested to increese it to {0} bytes. ZThe name of the site does not match the name on the certificate.  Do you want to continue? OThe name of the site, "{0}", does not match the name on the certificate, "{1}". %The new timestamping API is not found �The next-generation Java Plug-in option cannot be changed at this time because one or more browsers are running. Please close all browser windows before changing the next-generation Java Plug-in option. 8The parameters cannot be converted to the required types BThe password you entered is incorrect.  Certificate export failed. BThe password you entered is incorrect.  Certificate import failed. XThe publisher cannot be verified by a trusted source.  Code will be treated as unsigned. VThe publisher cannot be verified by a trusted source.  Optional package not installed. nThe required version of Java, {0} from {1}, is not the latest and may not contain the latest security updates. eThe required version of Java, {0}, is not the latest and may not contain the latest security updates. HThe security certificate has expired.  Code will be treated as unsigned. FThe security certificate has expired.  Optional package not installed. IThe security certificate is not valid.  Code will be treated as unsigned. GThe security certificate is not valid.  Optional package not installed. 6The selected certificates will be permanently removed. vThe specified directory does not exist. Please check the spelling or click the Change... button to choose a directory. HThe web site's certificate cannot be verified.  Do you want to continue? BThe web site's certificate has an error.  Do you want to continue? GThe web site's certificate has been verified.  Do you want to continue? �The {0} cache does not exist and cannot be created.  Check that the configuration is valid, and that you have permission to write to the configured cache location. PThere is already a shortcut for {0}. Would you like to create a shortcut anyway? ZThere was an error while executing the application.  Click "Details" for more information. ]This application has requested additional local disk space. Do you want to allow this action? TThis application is going to perform an insecure operation. Do you want to continue? YThis application will be run without the security restrictions normally provided by Java. ,This certificate does not have AIA extension ,This certificate does not have CRL extension !This certificate has been revoked 7This certificate has been successfully validated by CRL 8This certificate has been successfully validated by OCSP