� � � � #'<#9 /"0$3'8(5)6(7+<,?+?->,9)3)4.<.>,=,>,?*=1=[09X,5V$-N%F %D$)D'-?&+>#(=(.F,5P1C_4E^�/:U1/8U*3N$/N!(G7,3:YH`�<Qt?Sw6El:KpDTvNa�Si�_z�[z�Sl�HV�Me�Oi�Jb�>R�2Cj=O{0?p,8jG^�8Xt7[y:`�;^�7Xw5Vm6[n9_q!6(1L(/H)1I&.J(E&1R+9]&2N$-L*4P'=&<'?�)A'>$6#3,<f7Nw;R}E\�BX|2;`,6Z-4Y"*R$(J/:W)0I%);7KQ:MT<OV>RZ?S[�@T\@SZ@TZ@RX?SY?RY?S[�@T\Q>PZ%5E':I";F#9G(<T/Ea,CV0H^+@W,Ed*Dd)AY-AW0E`/I_)>S)=S-BY*BR)>I1H[A]Li�Pv�\��g��d��r��l~�j{�`�p��v��z�����v��|�����s��m��\�Vlt[l}o��w��w�����r��j��gx�_q�r��z��w��z�����r��bz�_lw[fo`p�r�������������������������������������������ȿ�Ŧ�������������������������0"3)?0;V=JiQ^�`n�`m�Yi�VW�XTz\Nv<Y�=]�<^�8W�5Oo4Pl4Tp9Yu9\s9]q9[u9^{8_�<a�js����o{�� � � � � � � � � � � � ��� � �� � � � ##5 0.!.%2'8(7+:,<->,>->2=1<.9-9-</@0D0F.C1=]1<[.:Z*4X$,N"'D%+I+2I',?$&<"&<(.F+6Q2D^4D^�0=VH(3P&0L"'B $>8.7De7Mm@TxH_�;Mu@PxFRxHU�M_�Oe�Sj�AI}:G~Ic�Jb�E[�2Ah)1Y2>r<P�FZ�Ne�9Yu:Zz<^�;`�7Vy3Rm2Rd2'0I,9R-5M*3N<&/N,:\'4Q"+H'/K'<&;#9&<)<(;#4"0"B2Ch6LtAXCW}6Ef0<^0;^+3])1S1>[-8U',I(-H6HP9MS:NT<PV?TY�@TZ@SZ@RZ@SZ@TZ�@SZ@AT[AU[?S[*:T'=S7E!5G'?W+GW,CX1J_,D\,Eb/Gc/E]4Kb0H^(?V)@U,AR.DT)@I#5A8RhBb�Fd�Rt�Y{�Zgphy�y��u��j~�b~�f��p��n��|�����w��������v��m��gtq��m��s��q��|��f��f}�r��l��������}��w��t��Z��j~����~��x��}����������������������������-��������������ƥ�����������������������������%( 0%0E0:RBNjSe�\l�br�RU�NDf\S{_Qyla}8V|2Qn1Lg1Og4Ul8Zv;]u<ax:a|:b�:`�=a}Km}Ml{������x��� � � � � � � � � � � � � ���� � � � V!/' ($-'1&2+9-9,9-=+;/:%:;5=1>1?/;2D2I/F2@`,5X1=]-9[-8[*1P*2N/:S*2F&(>$(:$):(/F'3M2B\.;V1?U.;T&1L%+C#'=&'@"</4Y=Pw3AeEW{BTx=Ks5=c<<nAFw;EkJZ�GR�5:o<N�If�Jf�?Qw)/Q#&QAT�Ld�H\�Lc�?aw?_{=\�<d�8W~1Ki0$*D0<V/7S-8Q!*G(0P,8Z)6S#+G#,G%9$8$5$3�&8$5!++$-J3Be@Ux?Qw9Gi8Gh1<_-9a1;_2@`1>_+4W)+I-1K5GM7IO9MS:NT<OT?RW@TX?TY?SW�?TY�?RY>;OU.C^'<M%=O%=U)DY'?Q-DY1H],C\-B_1H_5I]6Nd+@W#:M-C['@K)?G%4?):I3LeEe�Fk�@h�[��h��d}�u��j��l��^w�g~�y��k}�~������������r��x��l��s��v��v��n��r��g~gv�������������w��h��b��Ttxs��������|���������8��������������������������������������ƥ�����������������������������!(%4+0&%?% <*0 7``����}��y}�,HV/LY2T`8[h2Sj=_s?ew<dx<d~=a{Ccu^~yPs|Hj|Di|sx�s~�o��m��� � � � � � � � � � � � ��� � � � r#5#0$/'2(3(4)5