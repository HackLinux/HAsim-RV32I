USJXVKYYJYZJ[^M_bO`fQ_dS_dS]bP\\MXVLVVQX]R\cS_dR`dT`eTcdQc`Qe]Re[QaUM\SLVSOUPJSLHQKIQNGQTGQTGRRISUIQTISQHROFQMFNLDNJDJECICBIB@J?AK?BL?DM=DL>DK<BJ8BH3BI0@G/@H.?H,;E*9B'6>%5:28171708.7-6,3'1%/%,$*$*"* )'%%#" ###%'&&'%&&&&&$&'&%&%&&%%&''&%$#$&#$%%$#&%$###$" ""$$$##$$%$!#!"$&%'%'&(%'%(&)'*(+).+.,0/.0,2.3,4,5.706050314140424453535483=5B5I6Q6S2N.E*=-.".2$.4%06)28/6;39>6:B;;D><H?<J@?LA>MA>PB>QF?RIBSJCSMCUOGVOIWPIYTJYUKXUKVUKWSIXQJXQKYQMXNMXNLXRIXVJWZJV`KWbJXcIXdIZbH[_J]]M][Q\XQ[VP[WQ]YR]YR]YP]SLZIJUEJTDLUGOTNMQOJNIGMIEOKFPSKQ]OQ_PRYLTLLSALS<LR=KR=KQ<KP=LO=LO>OQBPSFORFMPGMRHJQJFSMGTRHUWHWYJYXK[[K[^L`cQehReiUcgU`eQ\`MZZMXYPU[PV^QYaPZ`R]`S_bTa`Ta]RaZQaVO]PMYNMVMLUKKSJGOJGMPGNRGOUIPXIPRHPOFPNFOMDMLCJFAIB?G@>G?>F=>G??H?AK=CJ=BH<@G9>E3>F0<F/?F.?F/<F,8A,6<)4;%2:27080:.9+6)2&2$.%,$)