                                   #Zisplomqvmlninmnimqmcilhhdddddhhhmdddddhdmmnkkggddqnkddggggg`egggghdd``a\``]\_\_]Y]\UPQTQUTSKOONOONOLHJH8888JKHHGPQ6888411H683                                                                                                       1_islgnqovqmqlqhlnmqphdjmndd_cdcgenlhlhhgmnqnnkgddmqmgggkng```degddmg`b]`___\]]\]YYTTQQU]SQNOLOQSSPOOHHHH888JKHHGSSOH68718GH993                                                                                                       %Wospdmlmyoqqqqhmhhisfdeqnhdhdchdhnmnhhmgmnqrngggcqvmgggnngd```eggghggbbaa`]Z[YX]YTTTRU_]NOKOOOPPOQOLLHHFH88HHHHKUPHHH8(1KQKHH3                                                                                                       !Uisoglqqvvqoqqninemsihcqnjdddcddhnnhgmmqsqqnknhhd{vgkggnnggggggfgmgeeb___\ZZZ]YYYZ]ZZZ]TQKKQSOOOOLQOHHH886H8HHKIQLHHH639ILKH6(                                                                                                       Jlwohqqiovovosqqqhelmhclehhdcdhdhnmhhnqvqqmmgknnmyqmnggkknngghnggfgebb\ae_]Z]ZY]Y]`cc]UQQRQTQOOLGHH8HH8888HHHHKPQH8H8318KKLH63                                                                                                       8dwshloqsoqyqqhiqmhisihnighhdldhhlimmqvqsqnnnghmq{nmggggnnnggmkfeggd`a]_``_]Y]Z\Z^d`^Z]XSSQSOLOLHH8H68858HHH8KNTNHH83"68HOLH76"                                                                                                        6dstmqqoqsoslmhnvsmisldhihhghhijhdisqmqmqqqqndghlvmggmgmnnnmkhge`eea\ea`e_`__]Y]Z]^]XXZTRQQSOOOKHH98H86868HHHKPNHH8368L8HLH766$                                                                                                        8iuuhovqspqsqnhlusnnpsjdqgmghghjhhlvnmgmnqnngdchmrngggmngmnqgdgd_deab\e`d`_e`]YZZ]ZXTRSXSRSUSLLHHHHLHHHH8HIH8QPIHH361JGHIH4(J$                                                                                                        Jdsxcqqvvnmsolnqvsqhqumdnmhhhhghhdivmggnqummkddnsnkggmgnmdqngdee```eb\`ee`ed`\]Y]]X]]TTUUQSOOLLHLLLHOOLHHLJ68PP87831LL9HL42((8"                                                                                                        Gdssgqlvuqesoqnqsonhlylhnnlmnnnjlgmugnnmqqknjddsvknggknnmdnrmggeeeef`Z`dedde`_]Z]]XTTUTUSQQOHLHOLLOKLLHHHL86ITL87838NH9LI662"8"                                                                                                        5_osglvqqlmqvlmvuljjiuignqmnsqjjdclqmrnkqqnkjdeoumnkgknmgmungggggeda`_`gd`_d`\\Y]^XY]SUTSOOKLOOOLRNKLKHHHL8HQPJ6731JN67HH326H6!                                                                                                        1`lnnpqllmnqvsqsxihdhomhnimi{sndfdqqmnnnqnmkfgivqqnkggnnmnqnfgkgggdb_`ee`_]__]YYZ]ZX]XSSROLHLQLOOOQKKKHHHH8JPPJ8433G86HH3(67I6"                                                                                                        Ughnnlnqmqlvvqouleceoighmqquqnhdhlsmmnqunnngmsvqnnngmnnmqqngkgggdae_`g`_`_`_]]ZYXYXTSSQOOLOHOKOKOOLH98HHHHPPNHH68668HH3269H76"                                                                                                        Pcgqqqqqnsqvsmmusjdcoihnmovzsnhhgqqqfnqrqrhhq|vnnnnngnnmnnmggegke_a``e``]e`]]]Z]XTTSQRQSOKLOLHLHLLHH76886GPPH6HHL69HL726HL72H"                                                                                                        Ncclssssnpoxvqluvlhiuqmmiou}vnnigmuqmqssnnnhlzsnnnnmmnnqngmnmgggeed`ee_]_`]_`]]XSSSSQSRQQOROOOHLLLHH81319NQJ869LL6HLH667H926H!                                                                                                         Ldclqqnnnqoyosqsulmoyqqmmquw{qlhniysmqsnnljel|ungnnnmnuunggnnngdeae`dge`da`]d]]]YUQQRSQSRQOLKHPHLH888581GQJH6HHJ98HF73666(2HH"                                                                                                         Pdhhsqqnglsylvssujcosquqmio{|qmnhqyvmmvnghdmpusggmunngnukdgkhknfdebege```_```]]]YVSRSTSRQQRKOOOKLH99816HNNH6HHH63H833$7762675"                               