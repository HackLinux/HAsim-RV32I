%�s��\>aT6d�%�宄bJ=�TOj�(��ۼ��e���a�� oD�S�΋
�����G�1��8��RMgt�m���3o���|!]��[��y(^�=_�\�y�k�>_9E�R�k����U��l�1���i��zŮԫ����Y��z��#!U�فb���9!�K7�a�^�B�x����� Ż4�M.و�(�E�e������ˋe-lhw
5���H�e.��s�}�0���9�x@�Z挝�Ĕ�2TY�7QXፚNs�3^�#T�e~�A��
n��vqϫ��l�%�-S���e���#	1�]����t��40��2���4�%_�b�Ҽ@�1[���D�,W�"jn	q3���N�c(��u�Pr����?��(6�;��]9�=��[{�;�9���4�/G�b��97�y��1��I��;�zGA.p���0�����q���?�8GWZፚ��8��]'Xፚ�^狜�\t�5X`$X��
?��4@��I�LK�|�.�@9�=�s$���7�{,�T�5Ⱦ�L�c�!�E��
��?.e�DG쫊�(_�Z��<�'���-}���z��0���nÒ���}��b��I��3U�S��4��Z�����Y挝[�Y���e���,�DF��P�A��
O�KJ�}�/�G8�<�r#���6�n仔�u��BA���4���"AF" �C��M0�~� �q�2Y?�t�4_�S��pwɭ��j�#�+}b���㺑�8�9l��	��B�$�D���2�$K�d��ܨ�2]�dW�b���䝶�{�]�V�����bfW��×�.^�ש]ፚ>]狜P[�Ո�'��2�`_�d��jF����s�3^�gN��h�b��K@&q�z��w�o���%��w��	1�'��2^>��\*'��2�d�D��(��Rq�>[�Ψ�=�������~*�Q�R��n����0�/�����s*���i8�BQ���nu ���薍�/���=U��B�s�<��e�%w}��1 ����ۭ�du���7�%@�Xx����Y挝+;��Z�P�etr���/ޘ��=\�<v�5XP�>���*��H�0z#d���M�����"I��Q��=��\N=:��Zn;>�$;׆��5�aL�c��{��=gU��B�3�?�$��ŰzW��#pl�v����/���%F�X��bS��D,�B�j7��)4P�b��17�T
��t�4_�.F�"jn	q3���N�c(��u�E��d.�e��b���
�y����I��y���<��\Ƅ��B��k���.٫F��u��{�zGA.p���0�Ѯ���Y��Y�T���|?��[	��y��(K���.M�1��9$@�S����w�4_q��FF��p7v��������r�����b��1��.��G�bs\�䯯�� �e4x���/ޔ/��=;���B��'F���vqϫ��l�%�-7��d�e���ө��Ó�/J^/�et�v�c�n"���c���/ކ3u�$U+�䞋�)�-_�#mop2���O�b/��r�s�����9�x@_)^挝[2��/��e�p��^�b�
��<D3��E�gS�cx�W�D�٭�p��|!Gv�C�����hX�}���EY�����?��\ E]����B[挝��s�2Yg%Z�����@0�~�i�ML�{�)�A>�:�t%���0�z�e^��V��;��.M�G�bs�6��y����~�x���;!���D��(D�by���o��1���i�������T��e?儍��4\ፚ��y�9��M�y��v�5XPD���e���7�y����LK�|�.�@9�=�s$���7��,�4�5�~��C@��Ev�0�c�v��H�d��>F��g�r�3^>6��E�$�N��a�$pz��0����ڪd���b��c���x����~�(�
�x����~<���x�C��D���n1ⅉ�⥵��������O�E�ֽ�K���A��a����
��t��=�����N��刮�����(���@������E���X�cx����{@F/w���1�֗�����LY㕈�⥒�2�u��4��	�BA��D��(��rs��v��p7�y�9t�����y+�V�U��o��鷭�S~�D6�E�����n�q�e4p������H��.M� F��+���C�B�F�e�����}F@)q��7��Q���r��x8���䣖�4(��B��3��yg�B�烌�.ٙp��0�E���*�`����O�E�ֽ�K���A���b��N���_�ש*<��[O�]狜���e�p��Ĕ�(K��r�3^��0�~��q���;Q��d��ŰzW��#pl�vb�A��d_�e�p�e6��ϼ��)v����'�du�a1��#�q��v��7�y��-�����y+�V�U��o��雭���^��W��o
�x��~�H�Z���*8��]�-v�5X�滍�/ު��=�,�B�pwɭ��j�#�+5��(�3�#H,��Dg��B���D�ė�2.�����~���剑�e�����>����O�E�ֽ�K���A�����*�?�C��SC�et�]��/ʛ��\���$ZፚN�p�3^�I�e~�,6�x����D�vqϫ��l�%�-���?��
�%I*�����X �du�<��(K���.�����:��N��Z~��p�3^0�GA��q0w��������pu��=��'?�~F	�;��Z8