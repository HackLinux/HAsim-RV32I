��F��.̛�.��U�x�H��$f����Pl�'5�5}�j��Y����S���\a.��#W�KYP(ŢX��E]N� �9�x��/�J��c��Ո��Xa�t��c�k
�̍b�j�SX���mJ,���;x���S^�#������Ԥ�H��Ё{XHg*Q���:-�٥^%n�����e���.8��/�dL�AI�4�yr�G`�z
>��(�n�3#y��ݬ(�}�$�	mQ)�X�8m18�>��,�܍L���\amѫ1V`!����*g��^ �^�{��+ƴ���`\��+8��J���̔BE>$\��#���HV�Yzl����M��ߒ����jyP`R�����R��㧡˦��l�w��+��0�z�'N�hI�R���q�e�`ct4�������g_ ��O�h���T�['[�T��` ��z�������-�iG�|�&DΜ��^6)k���=a^(����V)��0~��d`���1��������4��'�>�W&༅'�^|��u�w�����7���N���3�����H���&빽U.G���x���^��M`A.����v�	��qc	w����?�Z��$�\�6բ�O���}���r����D\�OT����m�d��=zӎ����o�c�!bЅ����&_���������P`�{���px~�4| �]��qU�4�s��x�~��?�;�R���.�H;n`&5戍�}d㠪Q��~�u�ĉ�+��e����ne���`x�B�b4�j���T��yz��b.1��6��,%X%�������H���o)@9�&.����6<���?�Ö��O��?_�ɜQkR,Tp��0��D�����h���"sN�@7e'�$���|�<A�)�\py3U�`o�������ǝG5l���
/ֱZ��f��/�����������Jx$�w2��+[��TE�'�'E��$6m�0̑i���i����(��'��ä���zK��i�ڕn�br�^�����n�FU�(b\��A���"��o�A���6���
u�~��9o�K���ЦQ����	Ix*p�_�,H��d���
�v�*�u��2C��0�M�of��hx������2|a�7��Ԙ� _#�@M��������n�^�g�P���M>�?��=���7�)��A���[dx�`��i��m��9c��n�^Z4d^{b"`+�U�,<�=]�RӶ����6�FFUq���ᩬ+��{B?�6���f�L�%�������MZ��V.�p�Z
|wFzT����ݮV7|�5Dٟ�>d���*�I$R��m�3����]��f��i��1�Oj�F��q?~��>���X����X���ItRm��%_:�(�G����	�ߘݭ��5��4g�8��[�y�s�E-��%�8��j* ;������6���On�]��wRya��MADԼv-����!E��*Em6����ѱp��F�{�H"u
���� ���a��mmC���_Z]JӐ\|�g'z =�8�bÍ��{D_��ph/��G���ZIife��۶���Ŏ��y���9_'�p��h�Qg��sD�4�0"s�Wܡ�O���h�ʡr�'���wm�ocu��{C|�Q����Q]�L��x���:	?D�^}0; ���~���|L�0�'n<o�,����Gy��T[����4l�(��x��ưs�v�d��~`or�p|��ۮ���q�L�^���j�|�?c\Jʕ|O�uP���zQ�n\�Z����U*���|�ڸ�:�4`��U^��W||�*:�t�2���6w��\)�c�]*�뼍PZ��PV���$!��d�(�G��9���ɾM��7eTBLs�h��(Ob��:������Jx�x��{�ǀ+�A�ssv�&�=D�q��V�r���'Cݿ,�(/�0p�,v�sSz̮cYm�p��qM��0��a���$��'$T_=a�ܞwJ�UϏsTH�Ө8C�gK��8!�y�@�8���}l��VMt*��L�]�p�U��+�Ŵ�e�_�����JM{��to��D~񟤓�|k���r5F��w^!##-���h�KGc�dG/��`�׺=��U�� B�,H!�!��.����b��hp�!� �.���Q�\G�֊Wg�o���t���=5��W5�k�zQ<(|z�Jy?)�@�]�R�<Ȅx<�O�軍��%9E�:�O�U#�_��Q{�*��%TBw�	��j�|����y����a':�0�����T����/��*j*ā�h�����o�N���_��\��p���}@E�.C�O�V�B5�n%F[�la��*���N_�� n�Mݾ� �!;��#��6N���}g��1n�'	j��I/��k4������%_�}-(\�����7��㺜d�w�� �7�����6�%� �_������p�������-�OL�������o��hT␆m*s��ɟ��Z%�u�a��������9���)AO��
��.A��Xx�j��8}O2�M&B�1�]O2jYc�����l�M�A�,q��&B��C%��n�%���ge|XP����&י��\�4�5�Y7��O��j?!zX+WК5J�W�A�5��T"/"V1��n_G��g��8���d�HN���a�Y��k��,�S��-����)� ��V��m)İS�JK[�M�G8	�{B~��QMQ1��B�BŜ�������\�"��ٹ�̑n��c������a��ƽ��sRڷ��{����.L�������d���b�E�����K=}���΅�`��Y�k��0�
���� �#����$!<Q�/r�1�HO�2��X1=t;D�KSf��d�.��=E�DR�f5*x�f��;	<$��=�[b��ϼ����=El{����^�;ݱ59�>�tSC�f�R;�<b�4_���Ef�����e�]�:�����"�� ��B8%�R�mUj4����b�"l
�
��m[f� kZa�����'�������l�2�z�p_�[B�}T�:D�݋z\d$�������+_栭�	`�Y���._j��hv<�6�}IG�����9��kQd`��Ma"�F�^ F2�`S�=D�o�[���>�9ŵBg���N(����z ad^׵BE�;�=�"�+<�fd��doZ���>/�S��\��5o��y}�U�;mꛃ����2�w��e9ߢ(T2���!��#~�F�9�T���k�>���w�Z�\��,B��o����EKWEq*^BU6�:J"iutpuc3onl3i{i{xnh3ejx3i{i{xn4~hswx2bkvtvi4d~jhyol~n3w~dj,/�acHȯ�y��%�~8��:hރZ_q+�{R�ՃT�2�|�Wԉ~}�$9Z��G�� ����{4�f��dTq��sיJ	p���5��Ăz�ڂPO��q�o�~=c٤`�j�`�g��De`��Eg�	���W^��8h�ԢHi�B%�7�D]�����Y�؟.�*���PF�����5��#��6����s\TU�D������
���b�_��)���b��;��Re�V�z��4�y��&���{���崠!q�b�MZ M$ϡ]�����8�����xcDl��5�^i�;ߍ�2�%#�P���"��
Ims�T�<<��5�����w9y4� "��^�����B�z��M�k#�~X��<?,N+��=79��[Z>�3o�&M���4Г��[^��y�dio�j��Me���e�CL��H����������˲d�A��|0O@�4��xJUx{�Mg���� ��~�7`�@�����ֆ`Rp�	���ڢ@'R�y.V2ó6�?a�iB�ٷ@eؕŎ��8�(��LX��F��Mz�79^�j|��g��蜴�0�+E��s�n'�ח1>̛�B�����6���~.�ʥt�,��R�@he�}K�W$�4t���a&\f��#R�NX��1Q$GU�/Ҫ��5x�N��U��b�M�"Q&��|I#7λ��~�,��I��)�~NR�"�&�,̷�'�_e��w�.x�������Et�6�cM�����`L��ο����0� ���[���\Pm!|�r�!K�|����.�~x������A�|(�Aw�iv�Z�>�t�d7�D,�� ��+�B�8����-oS*�=,]�_�Oa	� I���-�c\�jɼ���<���Z�ݱ�~/�2�	�SgC�UX�5��������a|��3����}���$uA���|�ιY@-��+�f4�V=(!V}1!��0y�S�}���%B�R*c�}NB������d<�V���\�k�|ђY�r9�HN`�n/����}�D����h�®s�('��}�4���|�̹AB'�`��c-�d���İR�%;�R�B�c�
���]����������T������p�к�&{�$�{0��?���Q��Y�u�G�����V�G���=�!��F9��do�Pf�[�`]�~q|�����\�c��Dl2�}�O=7bw�3�'��P�!q)�H)�����ن��}��}}m�0a'p���_i��j5�7�K)���J��'ޢA���]����Z�n٨�:@�f�/�ǋ�Nt5@߶`�U%`�b��O���`a���Mܙ�x�W�G��}e��̓%���l�mW����rըP�UK���]�XpT=>����~���%�2�b/�e����� �L}du_G�͹�;3�Z�bQǂ��JW��0LS��i6i��v�ͅT/0� �e��Y��8@Kż��mI�`|���$(#'#���(t�ڸ�ee��P��5�斾� $�DX�?3^��+Z=\#�E>��������S�5y+�ޢ�-,��c~d����=��UDb��$`~VF� ��圱�y���f�fh��=�\C����?~��Ҥ9�d.�b�#9�4ZӺ�h(�-=�mU������~�E9ɝٙ^������P-����
��$�`�������IY3�x