��##O�H��7��} �����"�)G1D9�AuJtSx\ee�mvvx.x�y�z|�|s}I}q|�zE{�zANO�##y�,����������
�e����j���w����u�Y�G�*������۟���'�<����y�,�A� �y�##��#_)"/�4W9�<�>0>;5�,�!FDM�
�X�%�]�5Γ���b�,�V�/�	%�-�54-�##?��j�!��߳���L�t���ZՁ���⻊�n�
������r��Ք;�D�s��ǆ/�8��� ��?�##���Ƒ��0�$�w�=��������義�b��շ����� � :�%�P��������������:����##� ¶�㲆L�A:GS��ǜ�7���:ޖ��iڀꀭ������x���-�7��c��p��##Y���.��� K 8 ��������}�u�y������ � b�:����������'�	������I���3=�Y�##�9�:�>�J��[�B�
I�6.�)&� ���o~�~X��js�j��g�6�� /��3f\��9##��}� r  ��7���f�����#���������*�����������P������D��������{�##>�5�)�!���S�'	��2X]���l��u.W�@A��"-8>##���1�+J&��M  ����������
�y���������e�`�(�+޼�7��A������##�{�w�"�G ����X�����������������������5
}��##��� ��������@�����7��V�
����\+�9�:A9:�;�=�>@>o;e5**��.��##�������������+�p�����E��N���^���_�3���
V
�	�����>W�##����K����j�����
R�3Y$�*T1�8	BvHLR~Y�b3buZ�Q_H�=)23%�N������##��]ܪ�z���"���H�d�c� wh�{^3� ��������������U�۩��צ���##��3�R��5���<�<��|������e�D�z���h�����&�����������g�����;���  \���  ��&  bx�      ��8          h      ��                      4          P                      `          |      ��          @      p��                                (                      8          T    p��$                  H��      �,h      ��	      @	|	�	      �	$
`
      �
�
      8t�������������������������������������������������������6�7�6�E �U����� M Q �_����� M P �^����� M Q �_����� M E ������������  ���?����������������������������������������������������������< �   � E ��a�����^���B �   � E ��a�����^���< �������e����x���b�	rL��	�a=����x��s�a�	rL��	���� �����u�1�� ~d� 7 ��L Z � � � ? - � F��� G ��= L � � � @ u� �������E�E�l�a��5���9�r�*������p����k�e��9���:�r� ��	�����I��D��ԟ�'����Y����+ه�2�O��Ԡ�'�����	��>�hϺʟ����	����������� 1�1��W������	����������� ���	0� ����
���K��� ��n�=����V���h�X�}�������� ��y�;��Z$�#V"m!�!�"�##��r��"�#:#�"G"�"�#$#�x��"Z$S����Y)�����E������k��������l,#�����E������j�����S�
�.f  0]�P$Vq  0^�Q$�
�.f  0]�P$Vq  0^�Q$�
�.f  0]�P$Vq  0^�Q$�
�.f  0]�P$Vq  0^�Q$�U,���J�����I�������F���-�6�
^��������a���n�S�����Y�L�UG7]/H*�(:+�/5�/�)�%�$�&+�0%5�-`)�'w*-/�4�/&)%g$�&�*^0G7��h��Ց�@�����ޘ΄�.�����>���3��4���ޘ΄�/��؁�9G�|��l�� �� ����7ވ�*:��"�T���V� �������7ވ�*9_�� `�� T?�H�
����{����\(�X��Z_���<����*�x�~���pޥ��ݑܒ���.����	�Y�bݼ�mް��3ݟ��k���h�C���m�0���c�:�p���N�r���M����S�/���d�:�p���N�k�  0]�P$Uq  0^�Q$ Vr    0]�P$Uq  0^�Q$ Vr    0]�P$Uq  0^�Q$ Vr    0]�P$Uq  0^�Q$ Vr    ������������       ��������������         u��?��F��T���B��"����?��F��T���B��"�u�_yI�l��a���������"yI�l��a�������������������������A�������C�������������������A�������C�����u�Q������\��*��ƌa��_�X��"=Tju�J8K�K�L�M�N�ODQ�R_�<����H�t�0�����R�Q�P|OcNVMWLjK�J�J`��烙���>�y�ǜ?���[@��wMDY��ޛ<���+���=�ȤM�`�6����c���r���x�
���T�����������i���$�����p���a���U���6��F���2�j��ߕޡݻ���'�Iڋ�$�J���y�-����ܖ�p�K�$������?����g�f���D�]�c�s��#��������������\���G���w����f�������"$^&y)-�0�4�8C<K?`B�E�H�J$J1H�EsC�@�=�:�7�4D1�-b*�&H#�",�	���B�q���+�6�?_IwS\�`�_�Y2S�K6C/:�0�&�`37���S�,�J�B�D�����R��,�ٰ�x�<�Y�����^�W��������������������J���Y����q���� �ߊ6��m��g�;�$� �,�G�l���΅�<�r���φ�S,S^S�S�SFT�T�T�T�T~T�S�R/R�Q�Q�Q�Q�Q�Q�Q�QR'RAR[RsR�RS4�3*3^2s1�0�/�.�.g.%/�0�2�4�5�5666�5�5�5W55�4�4V4#44��N� � � � � ����=d{��yeL.�����T'>'n'�'�(�)�*0,�-�/y2�6�;�?�ADB�B�BqBB�AA]@�?�><>�==T'������K r��	�vK��	�u A���h�N�b�����f���u� � |����q�m<2Y���~)x��+44.$	�tn7�	kg������_��H��_��,��%������s�+��t�O��5��k�C�"�����V�S�iHjvq]=��|J��o�����,֡���G���< 15���<�;����}�z�v�K�ϨڪD�㯏��k�M�o����/��ϗ�ֽٳ�"�����g��ۯ�!�tܲ��������ܔ�<���h�ۨ�:0�4[>�J�X.f�qlzn��uR]m=?�<
���6�c���~"�%:0\��  �                   6`          ~      ��                                                                              �$N          l      ��                                                                                                       �4t      ��(      \��      P�      �D      x��      ,l���h������m�����D����a�Q�I�-�p���g����|���.�����
�?�h�������  ����d�"��������� �)���Q�����D�����E�����8�����>�v�����    ��S�����9���Q���,ن܉�s��������3�>�@�7� �����]���-�B�  �?  <��j��
� $ ��[� ���\����,�    3 ��������o�I��������K����{�$���    �����$�r�1�$�*�4�?�Q�v �z��y    ������������!����-�Iံ�����5�)���U��6¦�tѻ٢�n����    ���f�R�t