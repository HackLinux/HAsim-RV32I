7F	#C�8㉯��!+�	tk���޺�ؾ�������_݂%��Z��݆�Eo�`���t�9�<j
N��u�%h�t��6 �����LӎaڻD�ގj��
�R��M����N�;c	�z�ܹ�\\��C}�g@�����Fby|�xx�$��}��2�a�C�}����L,[��g��U���[��.S�:҉��F8].�󼙄�>�|GͲ%���,��F���7R5�!j_�Z;��i��x��8t�}ߙ�A_�bJ���gf��s�������_�ٵC@�D7G��ܰ,$g��fÎ�>�,[/���ٴ��!����79���	��0�Q�,�e�Ĵ;���������@|fYM\�K����6ȝ��T�\R�F{,�d�~��p�5�Ǔ���X���x��:�;4'��&���A8#vD�5$��p��<� ��� O :��S58fw}�e���z�]�z[)I���.P� Ay萾�~i�lRpE0��)��Zz���R2���'�}R��K�w��t�}ŗb�J��Ѣ(��t�E^�(����Q�5�坿�'�*��x_�;���(�4t����m'�R��\�����%GZ/4�F��1ʄ��y��U��`��#~}���
\b�߰��#&I|����h1���5�MV� �>t���+����_�?d{�ol	�$��f�0i�²�B�����ke?^����"��������������/t��H� �$eE�޽7֋�+p�A�-�$Z9F��0��#}%ń@�~��_oL%��>Փ���<}�y2I�[�� Ȝv�%:Bh��H�7��<JA�B���w��1�(���a�Q��O���p=|�f�ZJEf���a����+�k#��Q��x�#�V��T���bt���~:��8^[�s����P����o����!���fǪ��pLC�7,�����a�ς��+�zy���d�^F��[��:���.�Z��܂��ʼB|�[`�w�&�R���@�p��0-H+��>��J�6���!��|���-�֌��;�@�QM�	�H�����
c{�����P:%��̋M��x���럞_t�e�m�V���ٖ�/�*���Q)�h�:JkM�Q��!F0�ؗCk�D�zBM��0I��w&�-�}E� �#C�~�f謦B��з2�>|ٙ������1�@k��X5�3u��=jX^��(�QVo����^�3���&��d}��25RKpZ)'������Sv��6Дcτ�&\Oh�VJ�	I���[���~sm��xՈ9��/����aW�E�=��c�����iu ��tp5�}����	R��H�wq����NDYs���	m�T��Z����Q�e:��{���r/]�S]~y��y@�qE)#�h(~��1�ޱÔ>Ѡ��+G��D�ĩ̱O��}8�Qwl���_K���u�ǇKx )�5��s`{qff�[a���N���Ew��c^�Ջ���2�������S���g2R�*�
1��T�|��jϷt2/D��'<��#���G�����+1L�c�[1!����o�G�H�64Pe�d~�)�-i�j�seY��xwq��o����mhR��fn��	|��;@�F1�T6-��R � �Ɗ&�Tg���?`
v@u�6{ ףB����V�U���:h���06j�ʘ��#��m��>�|�A�����sg���ڌ��[$� B/�f�8�:U�=���ާS��x���D��c-0�Lu��CKjDV>k��Sv�kk~�5Ǐ���&ى�μoS�ӽ��/�����73߱�����Â�����`�J8a�LM̵Ћ��\)Zc�~D�ݯ0A�YL7�K�p�B���82��_H�P��P�����o�%q�V/�ʹJ�W���7��/>����2���������o���!�WP�����C����2�����_l��a*j2���;�C�*�p-����2:y�v�l�O{{�t����S�h�߉
���3V0�U; ���Lx�M٣V�s�=C���R����+kE�#NXx+ad8E�6�ț�e+�ݴ��\�0�f-b�C�1a����ɳ�'�r��6��n���3vwȓ�t��=����4������҄fcL`�����꿩k���N�O������6�W��ΝVnQ������kX�澼ǁ�/`�%�<���XdORs�z�{LO��U�as�W�vc9G6�f��Z��R�H��j��+G�dN���x6ݺ��#l��lz?i��Y���︵t�0��m���ո���q��O�v.�AhVհGUA�cdʶ�Xnb�a��AHSHN���I���v6������M*������/��Dc��_�=Q=���Uu0���y�~�:G:2�X|�������������&U$-�4��l�ӭ~}�	8�=�9́2^�愰k��T�?޵�|�y�È�B=��X��*r����2�	����d� 7yIF�u���Q�Ɍqs'�N�Ĥ��{|M���y&sS�N�s���T�j�	U�jE2q*�u�`����^���A&/�Zeb=��bq>�)[(:Ƣ�ل{%l,h��mZ8��Cx�R�<p�T����O4;�gͼMNn�)v�x)�o��S`�W@
=	�^{
�i�S*J��h�҉o�(�d4r^���P���8V�X�e�]�f��<{Ts��4�t�}�MHj7�^�f�\�3;�wͺkF�Q�U}�ڱ`\V�Ыi���zu���؆��4�� 1��Y���T+4��J2�;�HrS�Ko���b}��[bꘙ��'q�5ͤkef��s���RhN0��&欐���i$���+��6Q���)4U;�=$��7�_�D�� �T#�x�AM�򩳌��B��<l��vCDb����AI�솕��{���`��3T���f��D�A���(~-[h(�	\B�3��&��"�S۔����Ȫ��i9jɸcs21��1��"�#�=�����xz~ �L5&��`7]��		��~8@���H&�;F��E����1����R�i���Z�%�I���`���AQ���J��U���š���)�K����cp���a�@/Т�Q�GJ����d�������E��ñ�=�T�c	L�#v���!��)
��d 3��˅���M�D�/%��j���h�d�e�Z��쁙)��
���aY��1��7T�W(���R��p�E�nx-������tEs�G���A�v�J|֧d��U��w
 +;�#�4�J����
��o��M�9S��[��2XVY�'p��"���k2!V�2�wZ# <Y�(;�@�$���������{k�jku:�n�]p%R�%��pk�sقH�s�_`�m����^Q��}��G���Q!A���,+��{��.q����U�*�SVf"�g�JSE�a�Ĩyү�?�Eu#RI%LzE8GA�Y:P�s�Ջ��F��0x����1�y6�'ogO:��7����[��b�G9��NX2��(�f�P�2ߎ�c[)Ͽ]��ǆ���[���K����W�?`a�
M�f������<&��''4C�@
M�x��+����(�D^U�$��[�UK�p?��T�9��Ð��~I�ܲF���g��q�b@W}I|��%�q�Cv9J��vG�;x��g�����d$�'&~��d/��W��d���le�i=�U�e��N���}2��M�3*f���Γz�U ��C���w��ޢ�����+�f��L�����&Z�&�0�4,5�����Y���זJ��B2Gz�[�0��v�K����Q�V��+����C�/*T�M��햩�{N,I鳨�t��UO@��<o����3�;E����x�=o)ů����^�m駮�Fy�_*�2��ŕ_���l�1̞/��A�Uh5=�ă�4@/n+Ë�R=&��:��_6 Ú5���}�[A���M�,<�Ef,V��}U�X�x8a9��AE�د�
B�X�\��
��˚_47�`W�K�Jlڧ�&�7[�7�k^�cjIL��Js,�m�;N����Y�s*����l�;�d�`}�l�޼w�t����W~�?|K�Â3���d�EA��eMQ�if�N�V�K�f;x�T�D���jٛ*��*�~�8A]vbQ֊�:����u��nX�6]X�6��a	����������E�8p�2*e㈐�[�e�gt��S�\�~�)s�G��� �>56���JrM2�sXp�>l��oݐ��3�P�!#�э�zQ�f0�1��a�!��5�{��>'r��E�)�9U���f{<�|o�lj�-�-4rzfj��A�e���#���|��b�Hr��#�2�w�������'W�3(7©Vp��ĵc��Ҁ7�̕�2u����t}�Lj�R���`�8���V�8��Ӛ��`������J��cWy�wlE��	���i��f:�g.��~�`+�.��τD�L��8��$OT�2[�8����0���ſ����{���	K��J�'&$��7�8�b#ČT랪��V����:5_�WE�E�5;W�0J��H�`����ޥ6��f��y�"���ʔ�]$s��9S� sN�}(�U�)�=9,���껈ʗZZfUq�i�L�?JtKER�F���u�[�.�~��}�uoJ��8��loxK��L& (�{�#^�a������!�y����{g���X.��BJ�����X�C*���[3�3��#�f����b��Ί����&O*�����+=�^r Ǿ��C��W����Vw~�,C,�#]1��;�l""ԇy�~�z�aV���,�p&�	�ML6Ǩ���Ai��h�\nw�´y��{��~����X���	����l^��
R`�z>���p,f1����r�*��|�ޙg2�����=�_L���y2K�6ٴ��.�}�um�x��=#�q�N���h�LH����^vĭ7sw��7�|\�S�D�Ye���T|x�}֏Z�Z(�"7�Z�	aO���-��h̀5n_vg8�n/���g�Jf���C�����(av���I�{��7�2��]{D݃��h�[��C�ы�İ�֭wB��wūv��~I�2o�)?�7�JӚ,� Z���W���0��+�4��X�*�p���.sK�p����~_�)ǖ���c�ԭ����k�n��dHtʾ�����#;�/��m�QX�F���'�����[/����W�)ac�7*�`���8e�T�O���d�nQ[�䃺fksڭ5M���*z���/��,�E�!���6�̓j����(���� �+��C�N�zd�>�׈�3 ��u_��}��s���m_ۙq�Y[*er-B�=M�V���*_uS��lfhm�W%T*�M't�{��L��t�:4e~���͕����<v�+���GA �?�wY�����,W>Eް��<��d�G���Nݼ`���'dϷ#`�o��IT��.��s����U_�2��(n��">�4J�_�LP�����Џ5�7�y�e�d?��h�GI3O�;SVF񽅥�B/�j�I�	�����'j�܏��j��n}�����������҆�V�d���/���`u��!���2V��+~L>�P���כ���v�������9GwM�v�4���S�����������0�����?���&L��$a�uQ��V^~��x��&�Bn��	7H! ��'!����N2N�&Igg���T���P!�����$H�WV��^ѹЬ\iV�^YI��x��`��������q�8��i?�q���~����nW��;C��HB2^	FQ�V#2� ݪ3I�qKΕLZA��ݑ�̨]e����:�V|.�qes~Bp������>��W~���Q�;ǿvZ�BCg����v�������J��j ��:{��~P�b�T��jmMM����v�����qrH1s�0���UDl�>�^CG��'��M��zbq%�d���w�����c_J��ߤQ�4Z�o���o��K
�eks�֏��͐F�q��4:���O���"R)��~o�ɕQ