���Ȝ�O�������ēgg����īj@j����dw����������ĸ�����ո�x��x@��x������Ԭxc��kj����ti�����psF-���Z������k&N������N7���������ƳgKu���ն�AAQa�����A		,)J�fS5q��������Ȼ~�9��������᪮꼦��xx������d���������ľ�������������xj�}���Ĥ�{�����������]NJs�޳���-''������Ъ����@00X��k,7��������᳇?@��᫆MQ������ГY0	 )$IE5CG��������~Dm%v�������ដ�ޓdgx��������w�������ξ�����ꮢii�����x@;�ć�d57?]����k]���rXd�٢t���_\�������puuk[E][jx] 0���������}a�ո�}=L������ĤXMja)	,RI$5<~�������O9l��ݘ�����uw���������z���Ԟ�������ԫ�����Ϣ��hh��ĸ�@[��[��N?@J��{kJoƓkj�Į�_w���١\?;��{����ԫ�����ĚAA����寸��j��ոjL|�ݻȹ�下jS�����Xw9v~�����2<��݌��ɗ�R���Ě����jX��峮�������ګ���������ʛI�Ḥ�raL����jax��Z*c��ՓCr������ٮ�j0SēJ�������Ȼ��ƚjAo�����ړtZQ���|)3�ݩ����]4o�����Ri7/Ob~b~���9<���q���Y7$��ޙ���ü���𧐞��������������������h��ĕjz���|�������x����Ć0r����tJ7;N0}}k����������������,��ᤫ���R��}oQ)T���O~�`�䧗�ɫ���iR�E/Dlm6T�y�6O%���Oq�֗?i�ϳ���ê����ד�����������ᶆ�������i��S����ӻ�⻻ֻ��L=����,xr@?1KK5S��A}xx����Ȼ�������ˆ0M��嫋}jJ5�x=)3bɩ��mDB2qm����Nj��̍�Ћ0Dml%6V9ǅ(�#���.9O������ų�š�����˓������������[4So��������o|�ȩ��ݨ�ݜ���=ck�����d 05J*K��c4}uu���ӻ�~��Ҝ��x4&[���ړj[u��}n��֩mO�O29~q���4z���w��a<lV9%��.^���((m�uJp����٤u������EMj���������Mj��������Ş�n��~~�`m~�q~�mq��LM�����xN@zSRsg[��j����ǘ�m���OT�c[[o���Զ�J{�գ���~2.~������z0���i����.`D.��%!H���..��s?w����Е\dxxa��j������������k���վ���Ą�an��`T�O�^V�eBm��j7���k0,�𤙧�����x����Ȩ�����OW�[[���˫xj@*�޳�Ȼ��D���~m��JJ��?���f�%^B2��H(���..��sRww����Z$Aa}���˶��������������Ԛj��Ԥny��2OmD�OO�O(O~ݶkk[A=����������d�~W(B2.���``�@@�ĸ��u�����g|����D22%HVO������gu�=5,�2`6!6ؘ.O����BB�swp����J$ Ld[[a������ד���冚���Ě}���˥���O��9<�HH�U(Dmȩ@&0��᫶�����g��bD#����vm�JJ�������᳼�g@����v.%<%B�?d���&?�x0/Qb`H%2�l#<��ɶe�٪dRg��ŦKJ*[��wI4*[�����ڸ���׫�����˕���ԥҘB�҅%<�e^�<.H��L�MY�����xx�rS��x���~D#����v�t?-������Ը���g*,��6(B:2<��?���Q4R=0�m(`V#(6�v%e������Ðj[z�x[A7@]��wwiiI[���������Y[������ՙ������ lҽO�BV�<.H�b�����x0Nj����0&Mj���OB##9Ը{g���F-�����ᤇ??t�kc������B<D%.���=4gXA0S�GeO(%6�������ސu�oa}o ,j��dh�������du����E}������˫��חӰ ��<~�DV�B#<B�bݩ��������姗aL|����O%.(9��ĐgZ��dIg�����|S74�gX�������B%9((֤����Nu�uMoy%mO669�6D��������]QE&0��0[���ww��Ţ��wII����j��������������D:l���BO�6%<.�9�~������⻩�����Ȼ�ݽ2.���Ħj,A���J����===$�>Zx���买926`�A���aAu�uA�bO6926�B�ѵ�����&&0A�xQ�������������ʛi�����������������66.^.^���BO�2%�.�DO~~���Ҝ�����ݻ~���H9������o��cR$z||��Y,p_��j��Ě�O!9.��A׸��u��S�O%^69%<�H��¸���&,7M[���̮z�����������ʛ����������������y�2O%Oe6v�H�B6�%O#�B�#2OG����TOq�����bO��.Db���ĕ��A?�n=n��}4?_���M}�ę��9BO�an������o0/�q.vO.2:%⥖���ż�R&,000Ax����Ф������������ʢ���j���������ӱL=yyO`�.��(�.6�B6%�<�%^B�ҽ�2(D`����<#y�`%m~���О��&������n[������zQ��Ĥj�֎&=�������[@�|(le(HDj��՞?��0@@,0Mj�������������������ʴ���@j��������ŐL4n��.O��B�.��B�!V(����2(l��ؠBy��(�����ٞ��I�����ӆ;x����AM���x[��΄j����x�;r�j+l^BB�zS[u��*EcM&;j�������������������෪���704���������|L�w��l(�l6�OO6�D�%6D.���v.2���Hll�B��Þ����Ja���������ګoj��a,j���R4AASQ4Q�jNQ=nḥeB(�;[��R@xrA70j������������������්���o7,@���������nn��w��^�l<ب� %<�9�%(O%���lH%(���҅%O~�Ťo�Ն ��������������a=S�Y �������}[jQ[x[AAjM[ճ�mq=�j@x�R;x��oSJ��������ē���������Ŋ�����0 �������յ�Yz��Iw�2lH��.:D<vT2.V%`����..vD��ҘHO����}M��a a������������� M	z����aMo�xja=0[��4E�a0A��Mcxu��*x�]k��jJ�������կrr���������������zz������ĵɹ�Li�hI���m���<b�~(�2TB<(���l�v.�2��ҽv`��®����Q�Ե�����������}4A;A		7м�A	jxjA ,���QE�[A��x��u��7X�������jS5>���������x���������˶���������������IIwwI�������Ը��� q<D%���26�(!�26�ǘB<���Զ��A=�������������}E���)	�Ƹ��z=AA;,a��xz��������ń4uc��Zg_����x{�׸�������������䥓������������ywiII��姵���������~2V.�ذ6��%6�`��V9���xa�oL��S&c�����ࢁ��jQ��A	*��ĸ��; AQA���į�����ի���� M����
-i_pRg��Đ�������������ӈ|����������ӱ|nwdI|�ֵY����jEE��~.^6e��l#��%��Ve��~Oq��Z4�Aa�7Y������ʊ������&-����aA[a��j�������ړAj��E7�ĺ�j7dF-
1Ii���꼪��������������Ӗ����������Կ|[z���ɥqn���Mz���L!m#%eO.��2v�H%V�����~~��s@x 0�A�������ii�����j),$7���ĆM�Y	a|z4jx�����ՇMo�[0j�ƓMSM0JŪRJ	F����s��������Ī������Җ|������ĳ��}�rS��yL)=���¶���ę�T!^O���Ol��#62B��`O�s_xx )�������τIY����jN$�᫓�Q}xLj���}���j	a��ExƕPX$$1"&FFFFF>"J�����¿����ĵ��騈|��˯���j[[Ez��yLz�ל������Զ�TyTOHl��vv��!!(.U�`9�̍s�[ Q} ,����ഴ�zd���ḓ}j>dվj}����a,,,,x��}���A��0@N]{N7$?�us�*gpw��Nx����֙����޳�����鹱��ڳ��c) E��������~�ȹ���פx#T��OeB������vD�2.!�ҌOm�ޮg7c�/o��������j=���Ĥ�����ģox�����x,[�x��ᓶ�ի�M&��/x@>@**?$I��*F�����������񙋳����������ݱ������x}z�����j�ƌ���b����}j2D�Ol#.O���Ǩv~޼ 2�#.���J}�M0j��į����M;˫}�������ԟ}LaaQ�ո��������A���dr��&*�Е@$0Rp">������������k�����������¥|n�����������aE��qeD2��ݵoM9D�x`l���Ǩ����%6.��9q���*EE o��իSQ�īaaj��,Y�ճ������Ķ�4)�ḯĸ������jX�ٳ���rN���E

&*'"F��ԧ��������夊����k������������xn|���}0;��`���цn99�LUl.B��Ǩ���gmOVO���˫x/0 ���oQz����}j��Qn����������o4a�ī������j�c?�������]'IF���ēa���������ϒ��xx�����xcjxxN��䵵�@&4��DG���Ե2Ga`Vm%(���դtg.(��Ԛ�jQ0o�Ջo�Ը���oa��aM��������˸�@,��������ċ�[R�����ه&*p�'"F���Ƥt]��Ħ�����?N]kx[���k[}�������§ӵ�m966H����m22c|ml(!e����k�%(%���aaQL�Ķ��˸�������xAax������ľ���M0o���������rS&"Z��us$&Skk���>*1w�sF'F�Ƥ���{u�tCg���J/@MNc������ޫ��䩻������O%B�vv�~��bB9��`v%B#%^H�ߤdS�9.2���[xz	��Ƥ�������ĆQx��������į����ԫ������whh��@j,	J��J$--?t����Á�is��ƕgguu����Ĭ�?/Z�k$[ľ������կ�q�������<2~�V^m`��v`e�zW`O22vOv�t?X�H92��֫���,,����ę������[Ax�}a[���ĸ���j����¸���ϛhhhIIcER��@RdRspK*-FFip������{gPN�����Ƭ//k5	4[@QS@x��������Ħ�`~bǰ���.%vO2��n~l(e^e�m^�K$?�DVBD��˓�o[0,����ˤ���ĸ�E00)z�aM��ڸ������ɱ�Ѷ���ʛhh8IJNw̕0jg1---J��������������K]��k7N	M����������������2`.~m��2%6O%l�~���n�l9el�ب��}7?�m�v���ē�[,,;����ē����ĚA)&aն����ԫ�����ӱ�������ʛhh8w,	7��g70""${�ļFh��������P5Z�x�߶����������������ա_�bV%vD�����B2e%O���ˆ��z0~`V^HU�����A)�eVq����c,, �����[@A���߆Lx�˙���˗|��������������ʛh8h�N��N[JJ*@���8����-8Fig7N]���ZCZ����ࢷ����変���O��������(B���}j�j;,=��:BO~�;)jį������Q )0�����[&4�����L,���䵗n|�����������ѱ����ෛ8h�&�ޕZ*k��YM���w�����'8i��**5C7@���tt�����������u����%(���帶�����O��oM@A,z����`%(���=[o[QMco��aS[ME50�����N4�����쵥����ɗ||��ԫ������¸�����󷛛�����N/$N���ɗ�ᮞ�����I_�áC]kk�{������������������ˋ5u��������Ā{�����նS, ������Ԗ6l��j4oxzc[Ac��Mz�oP50���A}�����������䶆�����ո������į���������x-����@7C*Z��ɖ���î�����pw��Ň{�������������������ᬚ�@>>��������į�������a))n=��[�������4ajr�xoaaxoM)SjE5/A��M�������������Ě��������������ĶaY������7?R�ڕ57N�CPj�YA���̮�����Z���ո��ĳ��������変����ϞX@Nts��ڿ����嶤��xZ��Ķ��A	,��}�j����a	4[}jQE[SNMEES;&&0 E;;������������᳓�ի�z���������ի]|��׭���Ru�KNZ��x��&4Y��pi����Ը������x��k��������������ʪz�Ԯs���ױ������s�����}����L	����j))Q�A	 QMAE@EE@00rj /5/C|�������⿸�����j, [�M���������ɱY0Pt�R7��i�K/]�����=4L��I��������â���kK�����{s��զ���Ϸ������p������nx���t���������Ƹ���Ķ��zA,; ,;;4 ,,& [}70&//��������Ը�}AA}0,o���������ė*?����{��8Ig*S��ӹɱ||��w���������hh��]k�{x��宪������ʞ����_�������}a}�������ĕ����ն��}����M,,=MA4 7/&	E�ĤQ;MS;/�ѵ������S&00j���������Z��ϐk�h8��]N��Y���Ԏ��w��������h���{{�Z*]������޳���ἳ�ڶg���������};j��������ڞ������Զ���ē0AEA)��t[E�����}���kS5S������n;]x�[L���������s"wϷ�{�h8�����x,����d|���������i��ڇPkZ�Ʀ������ĸ��ľ����������Ԥk@x����k���ĸ������Ĥ�����n����|}zg�������Ջoa����r/E���|,oxMS��}j�ḙ���ļ�RsϷF���ޢ8h���ֶ5���ă��������{��ޡ����NXZ����-$���tg�������u����ݧx[A|���ԇ���������ڙ�������������ߥY&4����֯��xM�����ݻ��ȥ0EE;;));j�������}x��������ծs��h������h��⻻�ٷhh�ո������]���������ī]}�Ħg[Pt��АKuu��������əxj������嫓������ĆMN�������������|YA|��y��Jtga�Ȼ���ȩ�Ȼ��ɧ}a;ALo��aa&7��������޼��_����⻹��������hhh�������{k��Ԧ������Ě�����$?&�ռ�>R�uk[����ӹɧ�����������׋�ԯ��]Q�������������ɗ����ɱ�u**����~�ݻ�~~��������cSA=L)	
@xx���������h�����һ��~b�`�߷88����{�����k{�ĕ{����ĸ�������N��]&*��x����ɱ��¶����������ն���}}������������ק����֗|n}u5n���TO�Ҩ�D9qbq~����jNS�aAj{�����Ȝ��ʢ_�ɻ�򰨌�qD�^��ʛh����{���㪐���{�ĸ��������xk�{7, u�k@A�Ě���������ⵙ�����ӵ����īԶ������������ն����ѓdNMM?X���m`O9�Ҩ�2O.DWm��L0}o}a5ZZ71u���⻜Ȱb�ʢ����~��~q~2%OVϛʛ��Ϧ��������ˇg�����ĸ��ͳ�xj70jcMMM7A����«������ӗ��Ե��������ĸ�����µ�����µ|�Ѷ��g\@E@jӻbb%9^<�Ҙ�BH9b9D��;j�*r�������ӻ�~ǽ`�����~y``ҠO2l(6vO�I8����ϳ��Û������x]�����������@&}a4	,����oJu�����ǈ�§�ӧ��䵵�������ڶ�����������}}]]gu�����D9(B2����(^D26�ݧ�0*�������ӻ��݌mǹׇ�y����TO�ɰ��Ǡ���"8h�������gh�����īj���ĳ������4	 LL	Lz���x?duj���ǹ��|������|�����������Ը����«}acQj���Ԍ��#B(���e%B2(.�ػ�**d����������ѱ�`B��}9`yDqyqTD��Ҩ��v���88h�������Ri�����������Ƹ�?I$$��j���n	)n|��ĕjJR7,,n�������ɵ��jnɧ��������ľ�����|ojSMx����u��^6(ǽlv<<2..6����0K���Ȼ������ʛ�l2^�~���93)GT�ǘe6l6l`�h8h��΋{��Xu��������ԋ����-8h8iR����}Ln����oA�dzuM7o���ԧ����|��z�|���������x}}��xj�}[a����J,	3n92.��ll2DB29����Pu�⻨���������imO2������y+GLb�ݹT2l(v�g�����͇{��������Ū��ޤ����I��h		��嶸�����a	M�и��������׵����jQz������ī�x����SMa[Ya������	Ac�.ؽv�HO26#6�ǰȚ�ŵ�m`�������hh�`Bl�ݗw��TqS������<~�J�����ᬇ�������꞊���ŕ��I*���,r�����Y,n�������co���a���0,o������ˤax�ո�[}�|a�Ɔ		A))S|q2��l�v.bGB<�Ҍǵ��Ҙ`V�����෷��~^(ցh8"�ߥ7{�g�����v�]��u��ո{�������ꤊ���̕�������  S�����yL0=n������˯A Y��x��AA�����ĤjA[��Ɠ����o�� )�A Ac�O`6ؽmO�9O32(B�ǌ����ǅ^9�������űχ���h8�{C*J�����kk*C{�˕�ʷ����������ЇM, @7x�)	 a�|���y=0��������寋A a�ΤX��,n;[z����A[}QM}���������	L������qbyBؽU%l(!%%#9��~����mBB����������{���88"�C*Z7�{����uN?x����Á�����������M&&@/&=)[}n���aL��ajE��ī|o��}�����ծd��;a�}a��jA))��)MMAY���=c,,S�������~`q%بeB%.(#+��yy+qݘH.~��љ���̞�>Kgi8888w{{��Z/7*�]PJ]ZC��ĸ���Ŋ����ᚕ���� 0MrY0E}���x����|)L����4j[AA4�������}x�мwu4}�����[ )�a4z  ��4Q;z���������|�n(�<<2#+i�ny3�vO6`���xgKC{�P5?��_Fi��𳉕k>/d�kk�xC*kĳ����������Ԥ�{���}[������Ƥ���x���|L�na,Q; j���oa���j4=��4$4���}�Ej�a)�"8���)Y)�о������������leOe2((3d����v~lH6`��J/*Z�57��x**���g���u�՞����k���g]�����ḫ��į���Գ����Q)})		a������ݱL,} A��A)Axzoj=�ϊY�ī�o[Ea��z�"���|�,A��4ASM��w�iJs���҅^2D63J����^�H9<O���*5�̊k���k7/x��\>?k���kZNJx��C$$��{��ĸ�����Ĥ�x����  =)	Lͳ�nYYy����a	)���aA[j����0[ŪIj�ų��Qo������II�z})Aa��ęQjokgwFiZRuj���9<%V2G4nye^6v��<���ᕡ�ഞ���������gk57k��kCJP5&N�k5]kx�������׆0&,a�ƶ j�4M��jd����ᤀj,4j������ո��4 QX����Ϫ[�ooj�ͭ��w�����Y,j�����wi��JduyO�H#.	AiGOO#q���T����ôʢ���ЋKg�ͬ����7*k��kJPxkJ[��k75��������[4&0;k���)	[��x4xj�������դ�xz�j��Ծ���LMg�dA [���٪u���a[aE�[$"$���4��A7dugw�����i$7��D��D+	AR36��]K{O����hhh���t*>ĕ]�����]{���k]xukxx���jN,7x�xN,Maxx������������ꮞ��udJ7$j��o��������awÞ&,��̼�ϼ��=AEA,M@?RI�ľ�=4o�du��gJd�����-}��y��|b= ==9B%9�᫐�|��󴢛���gr�{�����������ճ�{x��x��j@kN7N0&7}�����Ćx��w��ô�±��gRRR
k���������ِ= 4Ϟ&���������a[4)JS[�[a�������������??7,���³]L��������Չk`�����ug0�xP��KX�dk����ĳ���x��007 /&;���[;�==[@��ύIT�L=4&,&kxx�Jz��Ä?& 4̞$4w7R����ē�c, 	Kdu�����̳��oSz���I?���S,	,ws�{�Ћ>5����P{�v�����k/[uK>]��J0�k/P]u�����xd{�[;j[	&���5EMMax����YLTy�+	&@P/5}�dRX�u?E����dw�����ac;PN$>�����Þx}�Q;o�I�ڸ d�k07N]�]$J{\���������ĸxZ**����tNg/Cuk��*7]x���[xJ��zKg�������դXn��mD3=)?K*5g*
&��?JdR/C{��4$w��x� , Z���g���ٴR4}}M[z888w� 	@/7j���xkxC{k>*5{���׳�ճtuk�����Ԧ�d]rPu���&J@7c�x,S5>Jj��������Ȼ���[n�Ҙ&LQ)od7$

"$"dd/?	M;=)	,k����[$����R4�}���88h�hI��04*&�и�k�{�Z*/>P����t{�C$*������䳉g?������P	70N���j]�u����ֹ��ݖ����n�Җ=nx@,	)=Jc/*$$I-
	)			),[�����j��ρd��ī�Ih������]0&S@��x�и{��N]P?{]1Z����5*@���~qq~�ԕ>$���иC5*0][7&Qc L�������~b��bOb�����n��o4  ,A?*Mի5F'"$8III--
=�A,	&M������A�����ḋrx���������N@������į]���{j??//�����u1S���~qb`m���*@ֹ��7NA ]==nn���Ȝ�O2~me������na���nL=z����MM��z	$$Iiww���pK)���,;���ڸ��a,$g��АYE����ʢ���ڸ�}������ƚZk{{��ē��������ө�~m��ml~~�{7ө��]&, NuLy�*�ӨbGD%������=)j��|zY$��oo����$-"I��ρ'F_�-
  Lo4 ����ՙ���Ĭ�0>?X����������γ���Ƭ������J5Zg����Ȼ���Ȼ���~`DVOH6..2�{N�����{0*/] ,7]xZ4ǩ��|��O( �	&��Y4&8�Q	 Q|�-I"��4*"'�_1  a�����ך������Ĥ�kC*��������˸������@$]��d*/]���⻩��������yO2D<T�Z*�9T����kxj[x]kk{d|��~~����2!!H`�Rz4w��hY�x,		a=L*-�Fi�����Ю/)x�ḳ�����ڳ�����k5*$wg��o���������ĸ�r���P]�����⻩����~mmmHG9B<.<BHH��J5�D#~�dN�������N�ӻ�T�~H�H%2BDlv~�nuL34Y�������oa�Y

F"8hh8Y��I-_\Ax��Ĥ������嫫�����ľ�5*d�j;z������Շ������{��ݻ��ة�����~v�m���vl�vm��{PC?�~`�PX�7,���A	���ǌ�،���������ǥ*�L=z[[��£�������L
"h��ʛz�?& LSM���������Ḿ�������ڳ1
������ުp����u?]{J��Ȝ���������������������kg*&���`D��J��N	j��Mn����~���ذ��������zY��Rs��|n)	Q����A'''��w��ϷwŪ��I}���������������������*1�������_p�g*Ra�ݩmV������������Ǩ������*x���B#O���d7���/&�jj,nӰ��l%���ؠ������ǧ[�YF����ˆAM����--����ô���Ϫ$d�ô�_*	 	���������������������X���������_'F-'>���݌O2^�������vO.B�VBVO���x[z����~.`��Ԛ}ĳ�@[�j,Y�،96�������������J-Fg�j���������}>��--'�i8&"��	 �������������������u"F$�ӻ������>'-\ݻb�`V.9Vv�vlvl^%B:%%^v�������ݨ<O���£���˧��E0L����^2.BvO<Vvlv�����1"s��Z$J�������Su��$""IhI8hI44'F'  =j&$5����ԫ�g51$"?�Zɻ��~le����1'p��Ȼ�O�Ov.%2HVHBBB<.<O6.H%%29D~����ݘv6<�m�����Ȼ��oEj�Ȩ�Ұ66�l^vm|������>J����d>d����ZR�ώw���88I$?_8$ ,]@$77*7w�Ի����vm`q���j����Ȼ�b2�m�<..DB<<BHHH^VHl^%2.%9``q���O<(.m2b���ݩ������⻨���eOelqz��������77����Ğ"?����"FiR����w888L&R��A	=�o,	]1���О����өb~��v�v~��������Ȼ�~D(ǘ�`^B62%.2BOv�vv�eOHOVVODO���2�2B�2Dm���~~q������ǽ��vvO[���ݰ����a�Ր$ZF'8FFJ��I�����XIIhIh8w� &			M=&	&$u��������Ȼ�OGmmv��v��������ǰ�mO9Ǩ�v�vl2(<�����ve^����OO���V�(O�.2e���``O~~������˶�|yqGnx�����������$?�h'hs����=	dwg�Þ4X����h8hʄ�J	 $?d�����Ȼ����~W<^v��vO����ȩ��Ǩ~`eHVUO<<lvV^VV�v��^<��ee���l��،�(H�62V���em`mmm�����=		LL����%���į� Q��ê������?�j),{����Jp��838I��|	)Y��,n��м���іymqV.(D^: 99.9eV`OV`%%6<  v<���%H�(%(���.l%m^~����,	)��=,�b���n)t74a����������4?��oAii��zZF'��hh8i�, 	|��L|�����F$����mD�v^B %  :�B<.HVvl`l�%:%%V�^.%��؅�%9O#6���.�vm���� a|a	q�zM�nT3|��=Aa@}���������|�醁����8hhII�p''���h8zooa		|�,	����ύi7|��O��eVv�2:l!��6(HH<؅v��!%lB^�lm:6^el�#O.���<HOV(%.���69.�~����j�ո)	 x�g*�)	)q��na,��ę���������ꪁIIi8h��Ih��pK�ηh8n=�a	)��X"$��xZL��eB��l����v�����%9.%(V煅��2%v�����.VH2���BOlv2B���<O(����������a ;}���&�|�ߏ�4Q��,4;4}�����ś�hwIh�����Ť{��Ξhi�,��			*���u n��H���ؽ����v���2O<�2^�v�%��B<�ҽ��2Bl6#!2(���6e%l~%V���VnI����{}��Y������ZK�a|L)Ao��004,a�ԗ��w���ෛ�������oa���ń��aQ�a,		)||QLEj��Y;)��B2%l��v.�ذ(vǽ�.^V<6�V�HO2�؅VOllV^6.evOv<^%2%���v�BO~:2O���%I8�u��Y8I����_�����=Q�a& z����w����������=L�oL���zSa))MQn����Ƨ|=,E[j���BHlBB2266���Ұ�.2V^<^!e�%��и�|�%2#v�v��v(O2���<v�66<���n8h����wI883Ra˫J41���A��o��aa����I���������?	Y�	L��4 4=������ƫ�	 ����Ĩ�l6llV%DB<����ǰ(2l�V(l��n��7LV%#%(<O�^%���H�B6O����h88h�����߱ʷ388=|�Ԟ�"j�aa��==���ĸ��n���w���������4KJ �o	��R4	 	a�����a4) =���׻m9^BH�vVOvV.��%��ɿ�YymHH��3�7�<OV�l<vO ^(��酘b|�G6H�������n��������83��oJihhi"&�͸�������z��))������Ѥ��]p*,��a	a�Њ?		))�n)=�������ӻ`9#.^^B<l`^�ǘ%e��i88"?|q<Ҍq�xz��	a�q6BOlel!UB���L,;jrME����α��L J�������8��Y��ʴ�?*���)Q}ojoj���)a���ї�ѿs���xss_[��zQ���?4 	)	o�������`OO2����������22��whhhI齌��{��	L�����^H2vO<��		}�����zL�L	"	=���I��Ԥd���$��XA)Ao��ĸ�=}�����4���_���u����x=��J7Rdj�o�}= &����~DHVm�����v���Ұ.�΢��ʛ84@	 ��ԓ�j����) 	[��V<H�#lO��,&M��p�����|Y*?up>7AXd443hI���zJIs-7�&$u)	A�ęQ,�����)���_�������᫋u�Ъ&g��Ķ�M,j)	z���6el���Ұv������3bտ���豿Ε0$I��;g>���-=�l.(�2%vO�c7 AM;��'"8����-���ބw�8I$8'M44  Qĸ���վ�ڭ;c��g_������ć$J��w"�����ՙa,"hh8Ida�����y����xa���c@�����迣���]/ ? 5"z� IR7��#3[A Ax�j��I888I��Y"�����"���y8iůwIiN�IdA}��oY=,M=o����oS���uu������s-R��?$w��������a	=��88�������;&&4MxduIw��z0077$0>F'��Ԫ-&�%H^H��[)[z}���ʛ��ſ�Jdpp>?��F���ʷ��Ŏw���?I������a		,)Qca�˟����߶�}{�s>1N}������������M )A�LIwwI3	Y�����cSaa[uwhin�7J&		z*I$4/���F����"d�yv�9l6�ċjj}���������X*&c��K$?���������dœY�������4)=[x[,;[o����������M@J51@=������������n	 	Y	L��888I$Y����}|�������0@@&NE&		�����������1��b�!Too�xa��ĸ������a@����ꮐ���-����Iw�&IwdR��ݹ���o���Ɠ�x}˻���ݩ���䙆����������������,				�Y3IhI8I�������������ax�rM���?&4���������ոX���ߥxj}��������x����[a����ʴ������""p����""�j���Ǩ��ܸ����n)aS������~������׶����������}EaE04[}�|= =�4Iwh8h8>����������) �Ƴ���i84[a����R"*u�ոj*��Կ��������͸�[&=��홚���Ih�����iZż�h8T�|8w�λ�Ҝ�Ȼ����)
=E�~����m^ǻ��ⱗ��������͓]@M�o����ƫ�����o���hhhi
fr������j7E���u[���iI�],R�FL���gRwd|���������a[4��������Ihh����ˆ��R����wwѿwI����ݽ�������
;o�y����^.����俆j��Mz���ն�������a L��wIw���������u
)]}��ԫ�����Jn��ʣ�f4Ku��i-F-$����>���|������a�jo�������跛�����ˆ��d��������zI��~O�elVm����,0S��m����O(v�穜ߤu��?$����������j0��I88���׿���
c[j�ę�����II����N�����ϼ��K{���{\*��))A0|�nAQ}E=E��J������������َ������͞w��y9(O%.�Oq�˭���T6����H����يJ��dY����������jaaa��whh8n�=		|�=
E�MSQa���޿��8w����0gK��������*;�� 	C?��3),)a�ѥn|�j; 	$�����������Xxޜ�眩u��~VOH�`������O2����^���âi4?��7n�飫�����𙚸����ʷi��a,&0��}S/�ƆME=0Q���ӱ����  5z����X0,,7����|)y������ɾE)$-F''Id���*z�d����򜜌����~�v%Bl������~~O����O!v��9���R*?����񥇚�����o����������|u��KR|��,

}�帆x0   )AYA ;{14�������1{���|Y�������ɏ��F"�4 ,*��g���m~~���쌅��O6v�����m^6����6!~��OO�Ŋ[u����Ѹ�����a0j��z�������ľ�������oC
����ڬM	)cА>	zk�����*�Ŀ���}rS==��)o;  _F'wJ*44��i"��vV~9qyD��22e%(2b��^B.����`l��2b���u0x����Ḹ��4Ex��jo�����Ӛ��u�̿YRK
|����j;SE;��г�jwiI	,����́τZ����;3�TkE)	ks_Fsw��Xw��FR�(H`TmOO##�l�؅Bl�����l%B����lv��(D~��u4,,z��������EMo�˓[0j���zxtgJr�|R7\ |x SSC;�������َ,]zw�����1>���դQ����frS=�ޤXz��٪-Fid��s���dTmm~VHBv����HOevmUHv(vv���D%l��%Dm��������������[}���QE���nn��jz�¤w1I�K   	�a=AA[��r;��������	  Jk�śwh��J$Kg����L)���­�����|	XIii"-R?1�������q2O���.U<6<OH<ll���eH��2^2��s�AY�������������������|��||��¤R*"sK
	�ѥnn����};��K${��J	 	\]z�ŷ�i�ޮs">R&=��LY���ӵ����}a)R�J4]{g_p�t�ê�Y%6��e2vO(2%#vOe���^^��2m6�Σ[�aM��������������Ů���⹥�|������spFL��§|���|�����4$&A?P0	[�ww��٢--�4	n�+=�������ħ���AMd&Mx������t�����H2.6��v6�~vv(6vem���^%���%v~�ѣn��Y������ړ�j}�Ԣ�ww������ɵ�ɵ������ϒF
=y���A	Lo/�Û�iR���լ�r/N����pϢI-n3|ш=�����ɵ����| ;&,����������s1]NR��#B^���6.�ҽ�`^HBl���^%���#l��a��n�������AAAz���ʷ������ѵ���ӧn)|���_Y~�¶	 	 |�
���hI�������fCkg̼�Z7��wn��y==znn�µ�����jQ�aj����������F-ZRZ��.V<��v.l�l^VOO6v���V���%�yY��Y����������a[c�����������ɵ���ݥY,		n��>qy~��	 [E��;

��ʛ�I�� r��{P0�Օd��I	3ny|�z|=zԥ����o}�����œ������gRs�NgsiYe^��lB%6!(HeVv����B#���2�4X�}�����������Զ�������������ɵ���ac4	��Á=��ݓ0J{S�ݗ
0��٪��4	a�K  g�ud��83���ֿ|=)X������YQx���Íjjj}�ڼ���7N�di�lB��l.!2.^eU����V^��!~-'z����������������������޿||������}z?z���K
l��΀jx�|���C
n����ĕx0]�\>*$1����"3|����Ķ|@@N��zL�˸�����ʪudXx���êug�}dRiwD��`<bnn�O%^2O��lV^��6YZg$0���ڙ�������ī����������)	������߯�s7R���T���ԯ������J
4����ղ�k@�{kkPC-$��?i)�ӱw���Ճ5/@t7E�������ê��ů���ϴ��zccuwFd��|��ޙ�µ��2�U<^B��2}x�?���QMj[YaaQ4z��弼�����)3)=�������Ϫ7&����-T������n�x

�����Ю������k05t\���1����ɱ��w���g>0;@JEa��������ü�٤���ύdz�}o���uj=Jʴ��xJR����l%2V��2�o[7��|)S��a[M=0A�������=,n��[7Iw7J���[J���������L	 ͋
4AEo��KK�������fk���gg���Ե�豛��xFR?0ES[j�����������ԋ���ټwA�����œa,-i��ÞR?iw��6l��OچS;=�ո��x}��AjoSL�����L		���-$$?j��Y���I	y�����?0�,)n� �����c;���]g�᫱�ֿ�ş�tgP;)/o�����������ۙo���ުRX�������S[J$8�����sRgI*4D�����b�ԋ����ո��}���E���o���� ,a��-ajA0}�&w�dn����JZ@j�/0
&n|La���ڸQa��jA4��������Ĭ�sco;��嫞��X����cS��["4������𸳪FF�F"IR�u�ui4z���������������Ĥx�}����������Ϫ&$wwdM��F$?=j��M}�4	nn&Y��ӵ����0jQ|T���庋, ���ո�j,,��ޞ���ơ���c)�嫕��Ń��Ķ;E��) &R�����������Ad	d��������������������ՆAzA=���������ΣIXw��x��w?@}a˸���)XI=77n�����o];/,)&aY4@�ڬ�SS�͸����M��?Awz����י/)����������o0c�xd����ᮡ�ug���)		4Xz�;����Օ?M���Ƹ���	a������������ѣzw�����t[������[A��I&������&07&[��,Y4=�׶oo�ۭ������޳Y4�����������
�������޼;E;c��[����R'��L)	4wdw��������u &j�oLj�Ն=Qj�������������Ů�����ٞ�������ի�4 ��I	)�u���>0&���|AMRJZ���׶L/f�������Άj�����ݻ����ro������}0;S�Ю7;���'>sJ4=YIz��������x''* Ax��ojj��,)������������ʴ��׸������ĕo,��-n;[J?K1&*70**���|A@7�����=0c�ē�Y)&	q~����/*Sc;)/So��d����7x��>)z�ux[��Ķ�u��ok������Q		=��|	)aMA	    ����������������Q,o������a��7a�}]�R-�k/NNJt��Yj};@j����c0 M	&I4LA|ݘOD����>

;S��)4I����x��t?7����=rj@>?����������	@�׆)	)= 	)�����������׾�x���[a�ĸjj,x�����_'gN&@c7k��nYx�\$@���rE ?���|A4��e%2�~���}




o���=iw��M���_1��o=[;*t���zI��I4[[,Yn|-zz 	4XN,		*݌m~��������֗����ĚM0)Ķ&	0���x�K*&;�;�՗n���p*-*�����u��ӻ�YLY��~%�m���ӟ
S���=3����F"$)Q�����Q=�))N���i"IiIIw��|��n''*�o)Q=)=����)	�O22~��������|����Ć],|�z=������J0�{Z��||����$w�"������$z��ȩ��p&n���e%�H���ӻȥ 

0}��䗮����'?u���J44[�Ĥ�z4���wI���������ǖIp��aLSo��Ķ���j	�<(2��ҽ���֙������u&aē=Y�������{-$ JОФ���p�giϢ'I�ٴ�i�*Y�Ҝ�~��g4���Ol�������}
r�����h8_���Ydg��٢w�4J��ʢ����������Lw��T	E��[oj��SL4!%����(��ճ��ᦡg�����ĸ�E�ĕ\-$C���tsŴ��ZR��ʁ��ڼwh�d����```ǻ�Rq~D6v�������ݏE���7F_�_$���d������w�i�����������ʷ���~4��`+3=4��M,x�ċ�jy.%����~~������ЮZ$J�,A�Ƥ��&x�x>17*R������_�������"R��sw����И226����R?L�<6!6���Ȱ~��f
;���7$���ps���ϼ���II����������Ϣ����Y��3b��|��}}a�? ,��R�#^���~�������㊕��Aj����;Nx]Z?k>��Cg��__�ޮ��_""iig$Cg�v#���ɪsn�2(�����`G~�����zR�ٮ���٪���ż����&z���������ŷ�������vy����ո��Z	Y��%.���v�����ʷ�����zxcM�ī�ո�gg�޳5/�Պ_�Ϫ��F8Iip��6.vmm�����(��罨�Ob�;
������{t��Ԟ���J&,z߯[[)	Y�����������ӱ������鵗����7J1	��V%(���،D`�ȹ�hh�����az�}����ոg--���ku�K_���"8"wwi�4~%mOTq���9%6�������ݾ0��������o��ךu�Êzr[xr4Q��, o��۫����ԓd*w����T	|��Z�u- ���2.vH��بq��ݻ��������˸�����Ĥk--����]��_K�����F'8$��i�K=�`6v^<`~q�H%.2D%��^���vaaA/���������哞�����}xo4}�ĭ���}������p�_8F����^;}���̡sj�׌�.�2���ǅ~�ҩ���Ȼ���������ĸ�x5g��x�]5ճpF�����F��������O(O�D%9eD�%.2D~�L*�Ն =)�����������員�������,)��������ro������â�����|+Yzc}�����RX��O�(!�26�ǘB!B��D~~mb~�����������k@{�Օ�5��g���k��_w������ҩӻ^�<.<O2��V<.6H�a$7��aj	 7[�������t��xd���wIi�����㊞����u�����Ϯ�����w&n����Զ	T~2��%6�`��O(l�<~Vev�����������xZd���g7�Շ��А\��_8���������5���e2.`B���H22<�oAgduĸ�|d�/�����FMg�ϊIhi��)|����h8IIII8888&?����z������A4$�9��%��Ve��vOl�vD#������������ḕk]x��x5&����ĳ�{�����귷跷���>���96.lBv��eB|an|**wgX����?d�E�4R���\'$7R��iI�ʤj,��㴛��w�whiih8A����������4=Mod*|�Bv�H%V�����vvҠHO������������֋xg]���t/4��и������Ʋ��ŷ࢛���uJ;;�������b���On
$,[���dw��/[]u��_KP�uFiiw��Ϥ7	 �������෷ϴ�I"7d?"&&J��˸�����oS[a[Y�Vm��#62B��^D��H2922U�������]]���t/}�ᬕ��{��PfJ����ŷ�iF����uiiw�7J��êɌz?AM�Ъ���S;���̮����sFi���ʮ�E �����������٢g���ÞR*	 A�����Q[EA&��~l��!!(.U�^2V�%92BBH�񰌨�ǰ�Ԛ��{�g$��ᕚ�����C�����ԪFK��̢̼hhI*$Jwʴi7j4


-R*$������7j����މkZ����ê��u{;&4��������������������������ڧM��������v(2.!�؅B6eBHeOe���lvO�����՚]JC*-g��{]k���{1����ߕgKgd�������h�jA?��i*Xx07�ÞXg������Ej���٪*F�������ü�[;0�����޳a�������������JA���������乜~���Ǩv%    � %.���2vB������啋�t-��K//����g1R��īZ>KZg���������ęX��i-R��;a���ߤ�����ċ[���ʒ


-���ӫ������ę�j�]0;r0@@RRu����ī������}o������qB���Ǩ�v!:%ؽ.#e(e���%���e�Bm������զ>Fs-C�;�k5Z1�˕]1Kx��������ѯ߾�̢FIR��ո���������ɥ�u�[��Á����ҹ�E?pi�χ��kNS0c};@@d������˓]z��������k�x}j�|���Ǩ���%UBVO�瘅��Hve��v��v�6`������ճ{K'i��\����tK05uw��g\p����������������ii���������������z*$x��괁
����⹧N5RF�F7kxjx�˾�}����������|������ħ�[S07;A��񠆖�(%(��^%Uv2#eO��v^%HO������{Ck�����������@/��١K's����θ����������ު����}����ǩ�����$����F�������N/Ru����������������������������������j7/���3%��.O^2#mB�猘V2O.H�����ɫ�������ᮐ��ĸ�����s1g�������������������w���������������"Ԥ���F
��⻻�׸�X{���̐}������ӻ�����������������������M#2��BVv!<69VB��v��2O6lv������ӳp_�����g>-g�����u;N��Ȼ�������������ْ���ڌq����ݰ����������p_
��ǌ���������RJ���ݹ��������~������������⹹����c7	
~2��HOv%2..lB��V^H6^`����ݩɦp'Fϔ���-'K�__�Ϫkxr����Ҩ��ǩ��Ӝ�����г���~V����؜�ݻ������Ѝ�

L��`m���������>���bm�Oǽ���`��һBl`OBqv�����Ȼ��N*/�DH��^6^�.2<vV��^.O.B^O�����լuF'FsJ�Ğ���gF��Ϥ���ݨ�Ǩ�݌~Om�mm����Ը��D�����~~�����䵯sp'"u��HDm��ݻ����'"¨O(`.�e��O``��Dl��.<~��~�����ݵ&/7
Ѕ��؅~��<6#HvB�ؘm6H<O<D��ĳ���K-�����ՔK-F��p����mVVVO����ǽOH���������q<vBl�v``~�~�nAJF-�hR�߼_Z���ǌ����g

|(V%vB�ؘ<D2V�D��������`m~������M0@7@�e�罘���.%%9eB��lB62B(2�ث�����pI�����K$hFFt��2lv%2..9.~��������O.`Hl�BV~22`�AM��_�pF-��-F��ְbmm��u

�`�D�ؘ%O%��<l������  2����Ć
�9~�^92%O6eO��vOO%(!.�ɯ�ĸƳpi����{*77ZR�hF_g]�2�񠘨�����^�~mɸ���2H(v�.#vH������ЁI'_'FR���Tlm�ߕ'K�����ҨOl�.V��OBv!!(2~y����Lqm�H%((!.�e��v<2%6%%�Ѹ�Ƴ��_''i�ᔚ�u/x{sK��pFZ*&3�������Ǩ��ev~m����~2V.���.%V6�������ρ'hh�F"F__������g1''
Z���ҘHlvl��22v%�����Om~����n�H.22(%vB��lH%2(B.(�פ�����pi����Xk]��s'-�ggJJMy�l2<%2lHV�BB`O����m#V(���2%O%v~������ʛ'F��F_���ZZ\swg>'-*}��9%�vV��2%l6����ذ9.bm�����j
0)+2O(.lB�҅v%.(6(.��>s����Áps]  x���� ?pF����O#H!O2~���b.%^<���<9.~```��ݩη_>t�s���칈��s���ĉ�g

M��`mv(V��6%V2^�(%D9`�����-$*Y�2B%%V2��v�#6!#���gKp���''K* �x]tg�K�ôwLLy6�bB6H9e���~B%l^��V#(<2lDH9m�ǖ�̊?/{�����������������>\��|��l��2<62%B(^b�������i
�%.eH��l�v2.(�Ȼ�Z��tF]�0M��@7$M��Ϊ�_FI"I���J&4))G.O���U6%DB��.%B.eB<9V��~���/*������������������[A"�F'F_K*��%m��V~Ƶ�Z$&���F

*	%.OB��^Oe!%(�Ȩ����t>"*Z��xM����ī����Ԟ�_hFh��iI$i���l9%2���B6�(6~BH.^�O����N�����򶭭�������������êstN7]�������l^%B��{7   xg-''

TO9�҅O^.%.������k\-"Fg���������׿|�������Ţ����F"FiI&&*R��vHO%ؽ%..^�OB6v��9`m���R�����ڔK_\������Ò�������s�g&����穈m6W��NN5@/*@xjPC-"
?L^B�؅^v%(..%(��~�����F'�겉�����ֵ����wyi��������Ϟiw�����X*	&BOHe`l��O<l2.��B%<���O`T���pF���ͬ_F_�������ϴ��������̮�p>$o՚�ĳ�LL�x5@��������0��{0?K-

B.��l<6%6##%��Ka��������gCį|����������������������������"Vv�������ؽVl�2qn��[GmD��ִF���f��ps������������ϛ�����sZpK@�]*c������xx��������ᳳ���{g�R
)YQ*39%.~�1s������զZ||z����Կ�������ѥq������������JA��`e^V��vl��<�ɬgu?-ZY����R?��k��̼�����������㷁����-gt��{Nx��ĳ�ͯ��]�������Քr{k{����
sK!2~���FF�������ģ�n	n�IIu�������[0Az,LE[an�������������T<B��^Bll+�k{�����'$5x�ɤ1��\���F'_{��Ը����ٴ����uZg{]]��]xj�����5J]�������k5{������JKJRÁ���pF'����y��ֵ�n��IZ���{��g\ZJj;j}@E@o������ēNS��ĭ�������ȥ���Ju��ٞ/k����g���g'-t���55xĦ������gp���xNg��ĕ�N����x]���ĸ����]{��]�����٪F$����'F
F���n���ԶJ0�{*��&k�\KJ$J����d{���������{?��ī�������𤃞���������7����[�����'K���gZ�ƫZ>@CZ1u���k{�]N����{�ć>�Z7���5$�����Ἢ�FJ��R''���칗�����]*k/@J@kC*$*���������������ծ�Ԥ�x}��������R����������}����k�[�����_F��Pg��ո@5C{k$?5{�Ħ���J$5x���{@g��PZx?���>@������� 5u���֖|�����{57]{X]&����ᯗ�����������ă��txx�ծw��R����������������gt�,5>k������Օk�����5Cx��?]uk�����ƫ�r�Zd��ī�f5�{CZj]tX����J{����@/\'"J���x��n������k@?N]k00�@,zoc����nL�����ī����xgggR4�ts��dj������˸������ښ���5P������𦉤����ZZ���x{�����Ĭ�����kPN?5���j���kk*C �/��55����՚t\ "\���{\\��A�������ku]Zk70J0z�S40x�������¾����ċ���d0xu�dE�ի����������ո������5J]�]>{�峚�����g>{��������Z5Zu�ĸ���&����� *��k�5�f�CNg�@�t@/*7n�4���ͺ�a�; zx��Ƴ�����J˳a?�>�к��������Ĳ�74ͺ��&>�{P5,��P�xtjK*[7$-1*Yu}�==��µrY) 	a=���z�����C��̓�Zk�լK�������t�����8RǞJ*¯���j�@@ji"	)3;;���ˇ�;&������ͦ�ղh�����ަ�Лh�뺐������8��ٚ�@N\��--Z>F$3r��Ӝ��Q=�oG����������K˵�ꦒѼ�����՚�������$�w4��JF��F��$x��a�ӱ�Dǌ�����1�ھ��m~Ȩ�ƺ?J���厔����Δ{�z��ճ���ٛs�������/
p�����Rs�++C�o�yD�vv����ɩ�ܻ�vV6�VG҄F�������|�㊃��������]��S*�r�t��/
SK$��L)�ɥTA�,;= vl�ԥv���vT�vlll�<�<(�R8���ih�󹎱��p̔]����}��5�Jo1@�{{ޓsJ$P	�yJ��������L=Uq���Q=b=3H^elv�<�.%�_8�����ʿ���Ò��jJx�����u�\@ٲ�{��Z�,��,���l~�q�E|��=x� �	.66v�^�U+�Z��̐���wê���x{*kƦ��tQgJ��qrFg��pZuxXQ��7,�L2.#Blث���)) 	f{XS	H!�6͔ZR󮢋�Ჲ������z��_�޺�{p��XLkF���xz�[��ɻߵ	,mO����P{���/�j Co�O.��(�6��Z��̮�ж�ux�������гڼ��>s��"�Cu?��ӱ��)�����L.�q&�*��@y��k)	����|#�`:�D�Ѓ٢ʼ���������ᗂ��ƺ��F-�a=Ji��sA�MX鹹�,��UD�nn��ȋL5��F"�y���a�����E���y�ytjpق���������Ц�����p_14�n|î��Y��êdb��^H�a�Y��� �Q+i_���Q4�ͬ��k�?Y4@K��E���xk���ڔZ���׬k$��Ր�ju�k]���[��1�F"���l��YT	��C  A4iy�R*n)L�N[��}o@L���  N������]Pu��t@��p�>�g*��i�p1���8V��v��[7 �|7$=4$8�Y�I"�	_�sY/;;�CSo��a7Sɷi��㪚��޳��ZN-p����_�>����wO�na���X@JӞI�������w�n�L���[5S��`���Ĕ����t�����Jp$�F\����ʢ�snS���~<ӵ|o�j�|��4=?[J����˺�߆SococQ
;��2����	E���{P{��̾[@�k��Z����Z7��z[QΧv9��Q4ӯL��Rau�x�-4=��=������[|��i� 
 �)(��v�0�n/7��ޢ���X/�J/����r$��ZϕM��ty`2���p֯�wz�M�hd��j��������i8I�C9��v��}t7���hI�zZ)/uφg$;���K�к@*�b�j=�MM�1w���&x-i���z�������Ƣ���[
/�v�e6�)@�ڲ��k���A?Jp��x]��k����tt�0|�z���|jޫRX�«�w��ƺ@��x����ګ��q{N�ؘ�EX=���k tK/��{J����R��_?�xM�{S=�z�g��jM�|jI�ɭLS������Ջ�I������,�a;S۾�&=C|Mߔ�j�FI��t7�ÿ���J��$Z�t͝n[����uo�a�Q*	Lz=gu��ē���������º|�����}c��o������hh������w�微>'|ɡZ�M@굈ٙ䶇�꤆A�˫�4�44�������Ѯʙ������ы֎ʧ}a�j@&n�j���������ig��Z_�i1�70��|���������n�[��n�� �֓���֌�������}���M���ɗ���|���[x}�ݤ����������RZp���[n���k�����g���xa|��=aaEa����Ȍ`���ƃٿ�j������������ē�j��˳����}�[tï�IP��Ւ�];N�)[����S��Q����[4+FG����bB<���ބꆃ�����������ޢi���C��[?j�j��r���є7o|��꾧�n���}�ab㹩�[���p+q���##B��jX����uα����������h��xo�����=��Q�jZRSM}�������A���zZo=b�l`m�Ι��s�=l:^�!%D�B�z�̲ê�����ԧa�����|�ɩݨɩa|��j;71�Y}��~錖[A��g����62%m��Y����TV%�%(B�(�Xw�ゐ��a�����x���߯���~6~m�e�Y�j,�µ��x�`e�ǅyN���kj���v6`e�j�gzEVO(�%��6�pw��7Po�������ڭ�ԙ�vvlOv6�==;n�������(O��|?���Ԥ�AѠ#6%�X�4M=4<W(�!ƾ��d��MJ}_?���걙��ԙ��v�HlVl%mq��|���=z��.#��g�I���1n]���v6(��A0r#V.(�%`���jQ[E&�z�ʴ�p��|���ն��6q�Ol2O~b��ܩ��ɨ�#m�a�zX��=?i|��l(OQ��n�/�B6(�l㫪 &@���������ٹ����ǹ:(B��BO(O^%OȰ9V��<OO9����&zo�xL��j���`�&=���;�e6H��d0)4r�����������}�����nL~^�^.UBm%6��2�^�^̲�z$�������[�a��4)jn�j )�.V.}ku	>f&k���������÷�S4���Іz���ev2b.6��6l�e(v�z�=L������a)=���xoaYA{;�=m[j�	4n�X���헋���Ϯ��no���Ćui�6^�.6.V(%+�vlH��B����=�������Qj=a�L)L= a�a�����sa�4A)?�����������˵�����iXw���๧..#<�vB6#�O�Dv�[o|j,��٢���Q	dղo,=x�����x�A��,	
Is�՞������������֗uu��L��[�T2^O�U�BV猌�ZALG���p���[,[�r)==��ٚ 3]�/ �CJ7__Ri��ղ���ǈ����xc}�L|����.�U.ȅ�.2^�eł@|���Ã�麓k�����,L[Փ�}	�/,@?0R�*w�����������繹��[Q黗�����x<�^#U���9�X,Lc����j|o���ޥ}Y|���뫣=���@�a'?�����񓒴x�ѫ������co�(��n9ae!%ǰ�6(���, ��r���|� ����Տ@�����x&���L1-�ӄ�����sn{��f�x�ȶa�^eѩ2�m(!l◆.�f, ����}�j������a�߮��[-�R&n��Ji�?����kC�*)}�������6(vv��O�m2HvyJnD2���Mc�ͧ��o@an|լ���±��hh?)1�&[?>"s���t�}�r;|||����٣Vm��(.%%!O�kmV^��aal��Q,���n}ڇM��۵��������hho�4$$��h����C�Ђ{������TBv��mHvӓ�Y�^(.�aY}}��A;}��@���n��|±���ε��hLA�,X�|����pI�7C[}��������j��v�К�ߜ�4)}�����Mj}YroQ[/S�n������Ѷ��Եn���7?�[7@k�|�����࣫����߯���NZ����ѕ��Ι=qц=o|	C[EQ@0a //;�����͚�f4�������oxu*�wE��aA�i��Ѽ��u����Ѷ�ʷ�߄�륋�������=���o00=,&0�0,);����,G���ͦ1���hiE��ړ������h�r{[�����褄����a���啮��| |L=|}���}��E&f; S�N=˚��R���hw�Y���߯΍�j\��Z����������x[�������}������nA����o��ӻ��SS;=�Q;Y)r���С���卼�ҷh���짇����Ɔ��4��Z����ӵ}���ֶ�Χ������ɹ����5n�mǨW~���]QA|�ӻӴ��콩`~��h���ꕕ���պ���] �@a�����֫����߭�������љɱk@X�vDHؘ%<T~|a C�k��ȩ����~�~^.<n������惋����j&o,)��x�������������«����cj���.6��H%`�[|���ȹ�v�byym~ǰ��i8��チ��Ι��xd=*bJ	+��jXX|����Ć����Զ���xcn��t3!6�l%22l�|uب���yDҨ�9Lv�DHl�����������pi"���y�Yy�o������j���ц��oja�n+5TT��2H.m��Ψ`��ٛ�O~�Iyj��ߘ�j�����மR�n��ӈL ��ǲA��}�����aj��ֵ�cQomO�HO.(m��ǘD����Æ�8I31J���NZͺ������ )@	3r��|=Q�ѥ��Q���QaY�=�,4L==����T~6<L�T``O�z�x/phFn�|@*�]]N̦���ᶉ�o=oj|����L�==[=����[�z&z��;L�Y"�m=Y�j|��w��vH.A��vODғ&Cz&rr5߆Z���{t�M7��Ƴ�Ƴ�����z�nQ|�=j�Q4�&���|��Rw�3�rr�sipgve%(,YUO�b���ん���A�\X@nk&|���;,��	%n4|����xYx���nj@L�ㄋaML71�� zjdd���-Ay�T+4.B�zy󁛪J�{������{t��kEJMA}�������®dRS�����En=L��٥j)	Z�����x��sYM=n�L�{�͇|���X&jnnXu���z�0A?�A0Y;n��4�3*;�Z�tttZ*��= CA���XcQ|"h�	MAk�M@\&����{j���\k�,Ja�M&k����ɻ�n�3=,A/_*dN4	"qPa��,Y�?z��Fh��,)4A���k@KN��N*|����/��}@	5/&ELx�ǹ��q���nyC)�/""I$4	P���j��n�����r���x���[|��x��~m~�/��n)	LyJ��^v��La��)?�y���$-w�Ipy �쵵ѺE;$\��������X��5d�᩻���OH%(�;m��A@4=uY����#TL,=8y4	�aI�Lin$����߾���x/i�c�������{���Ș��qm`UV^|[a2�?LE�n3����WV���a3K�̭Ջ�
Fhi+"Qx����������C����[*S����ǽ��ҽ��n,j�.q�&�;kS���lǰ����ML�ǖ,|�$_�����?����������M"�ڻ�-_��b:~��v.H.6�����^v��Q|)��Blev���nRu4����/xx"*I8F �)�L;/$&-n���`��4?���`v.9H:O<OB(.`~Ș<Ob��}���vB`����n7��?ILw�$&�w88,i	T)5�����qvv~����Ө``�lO(%:���VmlO�vU`6��mm���ǹ~93�ۻ���R'FR�)w|�Jw�8w=	3&)n�ݹ�~V^26%bb�v^#6#6!##9eҨHe.e�UTl��)�YV��jY�����&�aM��Rw�-3�	T���,��l�B%�%H�#..62.l26��:H^�(Ol��=�3�43)��;Y�����瞊w8iI�1��wj			3K�,4�B����6�VD.�2OvB��UH.#�v6l%l�TTæ��4*�ǊwyaQ��04��Ǣ���ʹ�zӢRnL=)+f�onL;n�HBUB�H%�VHB2:lO��:9..:mvB2Ҡll6e�48l�8"l�Lw�LT0�=�Մ�����==3;�A&=���o,3��~e`eBB�H(�yTl2�y0B2B2OG��^qBvǴiw����II�nI$w��a���)q�ʿ��xX���	&)L����m6^vvv�U<�h8)����3��eV^H�3Qo�͆�	=T�iI���zX�ALr��4��|Ɗ��sz�A�[J	Y[ØBv�����T^�ôp)�nau�&�BU%^� ;�F?�~1wn44IIT_F*��n��a�����kx�"�뾧)ih43�Ұ�=A|]��===,3'==R)l.n4n|�_h�T&w�1i��ʎwy-wy�=4L��������>s|����;uIh3���LA���7 	4��Y�nyOT�n�����M=��\�@�﷯RnR��Lj�an����x[[������E))3_8F|�����=�x�u-	 ��jz�M4﹃��«Q|�x�Á���Ix�"�"3�����ֈS���v��ֳ���ΆE��n����΢�Mo�ٓa�43�w�	Jwn�dY����Lo����i����z�ů�"ㅘ���Env��:�ѻ��J��ƺچ4an8p�Y3�
 fr�˸4"��&Y��ӞJ�=);�)4��an;|������驲��<6m�ΜB��2���R�4�㺺ګ���Ê�J,d�;�[0LoqL  4=4L=�=���Ӌ,"$d)J��م����^O��O��.�v��4��֤��A�����£��Y)�Ɇ  Q�=3��i4&=|�amL=F?wJ�IL^Vm9vOeH�v6��6�em�4A�����a��4o�|xj��**AZ/0a0~���Yy���5	_��EL��}�� u�-Iw|�nO9.��(UUVD��2vBU~�L4��������ک���ȃJ_)҈�� ;�d�&	4)3���?_�qj��µ�=X4������!^�%mO(l��:�BH~�za���Y�â���ѹ˙T��W�LT
��I̱�S;��d�13�LQ|ũ��LEj��̯p?X�.e�%��^B��2�BB��|������������ɱ�|)�wl�=g� k�s� �CTw�i^�=)���|x�Ç���dgdDy�%H^��.�:H$K������������=T��Ӕ7��$�����{��aAu@	p{F�౱JQj=���Í��®zdiq�G��^B^e!~:Tg&�S�|LA����aLLL�n�u4΄���)���t���Pk�Z�й���K5A[�����ٯмd���x RʎR�B!~Bvj,�oL��an���=�4=�4�$T��?4�L= �̀E�\�����tS,�˺�ߝ��d4����uF_iwYRL��v�ӵ�˓�����в7�n�?J�|�LY���Q ==	��Lo�ˤ)n�����;0ȧ���Q�aA�ι���&����YL�߱�)n�����꣊��}���n ����	*;�4MJ��=a����A���������Q�|}�[JL&X�����"4==�nj�	��������n�ؿa�5n[R5 >@�xE7��=Q=��~�jr���t�tX�n|uj������;	=	������ެ��oL�;)��u$1;4��|��M	)��4�6^��o

;�aL��Y�w�)L,a�piRXY�I�)��	)6.���ۏ��{�L)���77��z���'�������&a�6.U�ֻ;
0�_=�MJ|Ò&ô����w|s����Q��l��لx���Q�>1Ő�w���_�����lD��&y6��Ȱf��5�Rz�����_�����÷�n�Daz|=J=y!�Ҍ��âɋ4|�n�\g��i��w'FR4T.~���#H�`~��Ã��ÎY�YaL�����񹩈Ǳ��X&�<l�~Ȟ������Զ?g�N�R��-8>pCnlT��.O�Ӡ�,����ڐ��xoM�=a���ސF?�)��Y�vU��O�~������ѬN��j&�p������Ҙm%V6D�.2#�&na)���⚯�̊�=Lҹ���������=Y|�)~^6#�O�<^eBv����ܲ]��k�Ʀ{���÷҆&�V(O��DD]Mp��@aMd��-��I�L�ٛ_iI8"	L㱗��L[7�`�<^酅v<^e���ӕ]��|ĳ��}��÷w�jd�z|��y*fՄ�C|ٍk�_�ʪ )������InRLJ=���aaǅ�%2^�<:.DHҌv�ݱ{]$�����*5�ՔR���ihAswM,
pJ���n���@?��ê{)j��̵������b�������^�G#�v^���ˤ1-R/��?>o�JP���ʮ��iR�Qa���ڭ��������k@c;Jx��������j;Ajؽ�O#.�^�26l��Be���xKp��٦NN��K�������䪁�������M��w��ӗ?pR���§��������ի�M=	�#e%(O��HBe���ъ�ĎZ����@��������ߪ������ɿM��i׽���Ӱ���������ݩ��a
.�:e.(^�v.:^��ȿ_Fo�K_������ǜ~���Ƴ�e�ǰ���ڲszvb�ӻ�R�~W^��e�lvOm�v���;/*L�ۅ�2.V�v%6<l¶�uY�ю*?i��<`6UVOO����DV��`U�MpR_�puӌ~�&
L2:`�<Be����y¹ Wq(.%^�^%!%V������AXZ�_J3͠�Ƚ�����%9�V:`���w"FFgzy�X$C���#6B�vUӽ�B~��;
E2!#V�e.2O�t���m�	&iY�B#:BV��B�e.Hl�ۿ_is�|u��Z?�O6B�e<%6#O���/)9%H�v(%!O�t�-'=�&)���4Yy46B�v.^�l.HBHؖ�/���������'1fQB�vO{0	�
+9�V2%B���K$dٓ�ڧ����i�i$"i�^�U.VBO�V�����t{��ߞ���s];�Ҩm3�NjS]�L@-D�W6.#H|�����S����������̊���U���vO�:y�^m�i���_������ôϡZ?�j��������Օ{}�
[%3�d?����Mn�����oay������Tv�lBq��-a�Mn{��_s���̴��ZJk�c���x[��Ƴ]�{��4>��") _����|AX�A|gJ]}[j����]�������z�� �A���-��5��kk/1�|u�M4�k�\7Q�k*��߮Y"�ꖦ��7X	Z*�곕����Ц�{�Ъs�������t M��w�{��rC�/R���xMZk}�j{j/Y�@��AP-��|z���kX]0N�oa�n��«њ�ga�n�������Ѧ�cd�{ޚ��]Δ��x����@��*�@7A nk[@?*&=a=��z=	f����{�tr���������"wL�aQJ&�-$)=�Ǘ=QL���˞��®��٫�ģ�I))o�j
"4��Xn9j�`���a�Ȍ`��p�����������}[4/n��57�L���,=e�|ba:vlle^I����ÎzM��Mgn0z��d43�cbBe�;�;3^Dlk�����������t�[4Xw��}���%m|C=L�))S�<~Um��ü�����˲�_=nX��Y̗byvn��)kI4�aTæ�}jYz=�z�Օ���X�1j�j�LuzI~��L4Y)4I�IL+s=Sk;L�a�ţ|�XM7$��)�Md̖m|��nzM=&mϮ��}S/
|e��=��k��[j\��[���n�`V�zY�n��1yu�굗�I&;)v�qC]ꛊ�L$��N�@��nL|Y�ju|�ni�|���岮|��y@�jzj�7�߇�@�J��a��|�n,LL��nݵ���|aa}�o)o��i�ѳ�zpNd�j�µ��|��L|nƻ�ЮվԆ��|}[|x��Ι��Z��z[o��z���Q=qЩV�Ӯ������ў�n�j��}��Y}���E��zn�~���TmH2��������§贆���n�aY����~j�u��!B���;OB:e��zL}�խ����Dl`oq��x�#~�d�za�62�nA0<(B`�jnA�w�їͺ�OeBmU�m�mB��M�=Y��OE�[;(:��A&o���༣��BOH6O2�D�^�|n���LQ�QnEYGLLaM�ѹ���Y�˃�B^D.�22�^�on�Ëa�==����|)��������z��̋6Gl�%V��Q,����a�n)|�==)E741��Ǯν��a�|��Tq%��a)���|a��a�֙Y�,&��Ä�����y�T|2vx.�Q�n}�����i&[4?R����A,=n�ٖ�e6<m|B�ay�;;�j�L������i?Y4n��w&aŗ��yv�~�M�|�,nQM E��ۺ�|����@�M|��̮����̪x±���=��,L==oL;}�) 0���d�i����٢�A�����󥆫������|�j~ތ�aQ  �۬�͈�i�㞥,�z�ӫ�ݸ���§nrm6�.G|,����y��lb���ӗƓY=L�}��ѧ�ߙ�n�L:�2H����wv�T�yy����ţwL�y����[�LL3�)G�bb(6y�v��d"�4Mzj���=A=b�aa|���L�nxLL|�wyO3qb~�znr�@�[k4�ˆo3)G��=�xnLz�L 4a|��XYyb|yʍoLr���A4oao�|=$|�LY��,n@nx?hG&goXN�n}�NLk;Qa����m&, $)ñ=@|�����g���yV9Q�AAy�#9GX4X3�$i?	G����z���[�����~TtTA0=Q����a4y|�)1�$Y3XnykA?��@1�lBlBH6~�V��||v.v��4d)zn$I$"3-=��vO2y�mH6!2.9V�UO~v�=(nH�=4i�,w|iIL4A4y�U%D!6D.:O<!.�D:my�Y=y�Y��֢_���43d�A|mUDv^`.Ua+29.#�lO�$�i3�$Tw|a�ʱn=T?=L�O��~yi)+nYsU2L)n|3*nInd31noǆ���xJ3E&ID�Ld�=)4n4O6wy�=dYY�nX�bAn�£[���QL3jI,j�z|n4�*�Jyìn����s�wL���)�~ǥ�ȋ�o��=T{rYY) LYaa=��=&�Lnǖ�Bv�vl�zYΥ|�o��|* 9/yaTwJ,�=a+?w?imD%v:`eelmX�⟱�ȫ�n*�)Es=LL�RTd��nAz�sTmDOlle^�����4�&�ao�QQ=i3�S�|����nX�6DlB^=n��[�|)L=�=4�nLP)�||u��z@��̬�j�YidD~��z��ю��|�)4�4 LTk��a|̈;��En�Xz&��&3noO��̗�|Ax*4M|,)�L)��YQ=�LJnL|uL4+� !����=a�Y*��di�X�~JU؈Sr?�n�dʮʨnTu,LB����o�uxn�F?3:�O`�E;����|jo����y|LL62�^l���{�4��J��T`9v6Mx)=�uj�Y��ii�z�jn�^v:e���{A��N���X�)R���zp�aA����yAӗn�2V(:�^߫>d�J�g��Ύ|��M�*��d�xo�ȧΧ�Qb9<�:~ꎄu���ǩǮ�����*����a������(ma=v::�(<ю$�M_u`lv��`lVOxs_Yyu)bWH�V6H��)#:�#6��IaMz3+6~OmB.e�Z����,[D~%#j)=+�..�}?����âdLY+O^BO~���u��٪]���x��{� &&3>��Au|znn�ц�~�y�4n4�d���nZzrj�nCLQ�Lu��j@)&|��Ķz[�����aj���jr��x}44LYA1=�a ������ó�4M�4zb[~�b~mY����|�nJ�ayLOQL3)(Wo�����djunw�ya4Jn3rLQ���[J�jnyy{zj=å|$=�o|�no�Y�nx|Yn����|E~4�s��z]|㙣aL�������x��xn��|�T~�=:V�|����v|y�O��YyTc3GoL����^OGO.v���=oabu&L���v9OmTL|�|||nL *�£��TyT|v0�|���?4M�YY|�~mb�AL=;�Qa�ju�����������|T~n=q��y���|=n�Ե|aT=H^��YYy�̆=nT��nL=jb=v�La�QxnT@Lx=�n)awY|c�bj)=|^a44*y�4�Y|ve`qaYl�LaY?I@~BGH.:6mV�3Qq[zww)=yTly3L+6Tn=iLLTʪa434dnn,)YT��nn�n`�����a,LL==nL=YyOByln�̿�L==EL=Lz���DT^^a��nYL=n)=n��a�|xAnTwy,��on4z?LTLTQanu�T=A.���xLpYD`3Tk�z|�nynOD:��\n���4��Y�|���T G9H�gz���~yX�Abm�9LUHYYLy=OOD���LTyz�n;*�YA|��|�|a��j| ����ڴ�ښ����Κ��|�����w��uҿ���\ߵt���νX̵z׭u���ߥWƩtޙs���ΥX©_��q��������R��F��^�����n�����_���эT�����Q�����WЈ:�����\��J����R��:�����B��J��;�����u��L��9�����B�hN��z�����B��{��O�}0�{9�|9�{B�{{�}0�{s�|9�l*�{k{{s�g@�s5�s(�sH�s9�s1{ss�s(�s9�k-�s1}qdssssskssc�k1�k>�k)�k1�k!�k)skk�`skc�k4rkZ�k)�c,kkc�k!�c!�K)�W)�c)�c!kcclcZ_6{c)�ZkcQ{c!�Y�\�Z!c_Z�Q&{Z!lYN}W){ZsX/sZ!cYO�RrZ�G{T{RN!ZVRpR!sRcS8qR~IkRWRJ~GsJcRsJcREkJoJkJ\I>gH%RJJcJcJ�.RI=aKoBZKJJBnB�6cBcBWC%cBYBJB>NB1n9
ZBZBRBc9\9B>9U7$^9 Z9o.R9R9"
R9J6(R9 B9(]1>91J9V1W1 R1J3]) J1X)
J1 ;0,<1!@1oB1R) A1 J)Y!J) C)1-)<(!B)B) 9)9)-*!J! 9) 1- 1)1'B! ;!Y9! 1!F 1!1! )!%!B	(#9 &! +1 +@ ) !1 ! ) $!  '  	       xeno_sup3 a     @   �   (   (   ((  (*  0���n~��������ʸ��Ҿ�Ҿ���һ���δ�������Ҹ���Ҹ�����ssʸ���@@S@ f���Ҹv��������������Ҹҝ�������������Ҹ���ᇇ�Ҹ���ʸ���Շ0#9SS���n`n���Ҹ�Ҹ����Ҩ�Ҹר�����Δ�������nn�Ҹ�������������9 ,9f��ҟ�����ҟ���Ҩ�n�����������΅$y��������筸�ҭ�����������#0:~�����ҭ��ҸssϨ�n����Ҹ�����T>���������ʇ��NHHH\���ʸS 290n���������Ҹ���г����������������ɳ�w�D"7Q=GQ f#-#0:=^kIDNHHz��uu\lh}||�������l$b���|]AD7'3Fg;    S0#-@!%/&3&$*AMee����ֽ�T?j���]**?b�������ޗ/ -@0-L:PPPQp\F&&3Tr�������������$)������������������۵=!-:0-#0@K 0SB.i������������������������ڋT��������������������ʢ��~Sf@#	0ff����������������������������ޫ������������������縸�Ҹ��SS02#`���Ҹ���Ҹ�������������������ƅj������������������ҍs�����n#fSL0n��һǸ���������������������ٛe���ֳ����ǟ���ҟ�n�������ҟS- @n�Ḱ���nn�Ҹ~���绸�Ҹ���ҽ���e���ɜ��҇��縸�����ҕ`n��##�ҟ��~������Ҹ��Ҹ�����ʸ�����R*���ٯ�縸���⇇�Ҹ��Ұ��s�,f��ʸ��fEiwf���Ҹ������Ҹ�����Άy�������nU������ʸҸ��縟C6SLf���zQD/'14F\���������������ι�������޹���pz�IwPB�n`��#@@+:=//DD''A\h��������ˮ��֧���eb�����\D/"";///I.# S@K-#2^��������r>11>F\}���ўr��ַ���l>$)>DT\r�r�lF'00K9 Q������������޽�ll�˹�R��ޣ������l8�������Я�kLLU00:@@0#.�����������������>*����^����ȹ���ֽpw������������SSS9#0@S������������������pr�ַ����k�ӷ�������������������������S #0S�������n������������������C��������������ƫ�������������S#@S�ʇ�ջf~��zzz����޽������������������������ƌ��҇�~d�����f@SS�P-/ugVA4AAA3;T��Ά��������޽������������~��������һҸ���.U�90@S,,:h\F;DYTFTV\Y\by��������������������s�����j�����Ң�mD,n0@S:-;��������Mj����������Ư��ջ�����������j����gu�iQ/#9������������Ƌp����������������⻵����������juNgrNI7@@S���������������������=!!!!!!!cr������T1;FF3/+n��n�������������������Ɗaaq_aqqqiQqqi=//������>$b�zwi�U0n�Ǉ��~o~��������������OOOJQOOxq{O��{aXQq�����ΣRr����縟SnS:@�f��fo�����巽������鼈Oxxq{{{{{�aOXOOXO{X�����ߒp������Ұnn+ 05������������*����ռ���_Oqa_xx_OOOa��{Oq{qO{q���ٛj^+o������+C~�%%Dm\\\\�ѹ$���ܓ�����J_a_xx_x�x_x��J���Oxo����j)p%������LS�P !&&3NIFh�e)���ܑ���xvJvvJZJ_x��vJJJUJJOJxo����DzPQ�����#C�//D\\����YT8����������Zv�v��s���Z����vUUO�������p���������(U�Gc������V�����羍ss�s�����s�������UBkp���������ƯkPP���@ 2Sno�͵������֫������ݾ����������������������������ޫӯ7 nK0@�����ͫ����������������������������������������꽣�ɒU0  0: @����������������������������������������������b��ٵ~@@ S#0~�ʸ����1���������������������������������������8T��rk`LSL###:,^gFF\�ٛ$������������������o�������������������T);DNnn�@@@@L'4ȹMM��������Ң��O��=q�Q�����������ƫ޹����֣I7Y��`��S#@LEINgNY}le���ʸ���ooki!�Q!q�!��q!�������������ƒwi[i�����SSG�����r3*e��������������k!���������������������ʵ�������n#:=w������ֹr$y������������������������������≢�ʢ�������ɵո:@@�����闧޽Y������䳵���������������������͉��縉�������ւ�SKn�����z��ޅ������ޯ��������������������������ո�w������zi
0@�ǭ�ҵ��ޛ�������ʚ�������������ʢ����Ң�����Ҹ����֌��=:f@S@Sok�\h��ֽ��������������������������Co����������T�νf-@S0##SP\F\��������������������������������������������х)��^####@0##@~^����Σ���񟕕�������������������������������˴��lG --0:0##f������Ȯe8����ʇ�n�������������Ǹ������Ƕ���������ѹ1G##-9@0�����֌r�l*e����޽̽����������������������ϸ��������ꋣf:00(n�������Y1>V}��������퇸���������퇸���������ܕ�����t5#	@v��һ�����j�����������܇����������܍����������Շ������ނ05#5		n���k����ތ�����������ܝ����������ە�������ջ���������T֫iC55	#ҟU/���ƺ���������������������퇸��������镶�����$�֚S5JCf!/��ѷY������������������������������핶�����*��##,50A��х7������������҇����������ׇ����������σ������$M�K
5# %F����1����������ܼט����������ϝ����������ϥ����ˆ^,#0	,:@#-I����y$������������ܟ��������ܝ����������ӷ�����*$$B55009@LG�zrruy8����������������������������������������lM>r^S6s0@SS0i������������������������������������������������������o��-@00o��f������������������矸���������睸������������������ʸn#Sf~ʸn������������������ܟ����������ҟ����������ҝ�������֟�C ns��v�����٣������������矸���������睶���������ݝ����p�ޫ��@#CS���SK����j������������Ҹ����������Ҷ����������ҝ����)�ƚ�S#@SSU�ҟ����R�������������������������������������������S#0,#-B~�����yr��ӣ�����wt���������Ŷ�������������ll���D��S-#S# #..=kr�֣R��}���ֽ��������������Ŷ����ʰ�����eTTleY!-00#:C./34V���1?��������ã�Ǹ�������ŸŶ���ǰ����ι���Y@@9C@I�����$8��������������ҟ���������Ǒ���������Ά>TVFNgK9@KS@02Ip������l*b��������������ҟ���~��������������֞�������n:000Lo��i������ֽ�������һ������ҟ��PPO������������������ͳ��@@#S�����җ��������������������Ҩ��B�������������������ޯ��͉#+0#���dS������������������������������璌��������������޳���#-@L���ǟ��z������������ͻ�q=��o���������������������ͳ�����## 0@�ʸ��n-Qz����������ͻ�XQQ�t���������Ə�����������ƫ�US5K
0CU����K0f�z�����������͠����w�������͉ʞ��ι����j��޳��Ҹ�S###0@Ln�ʸnnwm����ӛ�������޳�⿒���q;X����ή����ѹb���ڳ����L0,9@n��S�������w�������iPʿ���"=Q���ٹ���l*1�ίg;0#:.G^���u���νj?�����oOf�ʣ���/�������ў1$l�r70:##0@SP�F3"����}18�������P�����=���6����by�ѹ�gN..=:0#@@@SCSL�c7""7NYFVYh��Y��������͒��������Փ����ֽ�����������ZL@KS95LU~������������������Ӓ�����֡��ջ�������������������S@@@L0Uo���������ճƯ���������귅�����ɔ}�����������������������:0:@-Sn���������͵������腽���宆�����ޞV����ߣ���Ư����ʟ�����#0 #^������ҵ������օ��ֹ�M������T���֋��������Ұ����� -0@#/BP~������wz����pT88e�������T>��jD��������ҸʇL-0#@BSPPP�o�������cz�����Y*j�����ޅ$'>1j�������ʰi^. 0::5U����f~��������kc�����e>7Rl����l))�����յkQgN/:.0-0+-@#@n~PP��i���������i������l