ddd<1Uiz}��}}}�����nd�����������������vv��}tiddq}�������d*(LU<}������YD<%'O��������`q�vv���������}}�����������������dWLLEObLUUWdU1<UiU}vk}vv~����n}��r�������������}�������}v���������ibindL�������\1<?*%2:O}����q��v���������znz}�����������������}idWOdidWLWddWLWU\iiiifk�}}��sn��r�������������������������������}WRi�������ngWF<1?*'*Odv}k������������zii}�������������������}pdWdWUU?LUddOddvd??Wikv}}��}n������������������������iUv������fEL}������zR\WLL?6828OWd?-Oi������������niivk}}��������������}}}kiO?<<<<<<?8Li8O?<?Udkf}����ni�s���������}������������dd�������v`}��������}p}fdbL68OL% 8d�������������}LLWLF\p�������������v����]86??6*%%*8<8OfO6?Wfd�����n^gMn�������}Wv��������������v}pk}������������}iz}}}L%?dkfdVO8Ed������������rU?<*Wis�����������������qOL8**L88661L8%8Odf��i��uUU^������^F?i�}UU}�}������nWppu�����}��������}U?bUUidd]VlOLUb}}vv���������U"OLddFi������������������v]G?OOL8%%%28]]fvpiv}�\W}��zK7???U}zD<DDU^\WdWLLnnz�������}q���n����oOdv}dL%%LdWbigi}iU]��������WVvqdL8i������������������vfvqqvd?%%88%'0%G`kv��nnnULz�\HS\iib<UD//*%-L]`G4Giin\n�������i��i�����qv��L %*6<Wti\Ugizp�s������}odv�d2q������������������v������}]2EL88'68fv}��UUUFi�����}}�}ddiD***88G.2'?q}np������v]Oiz�����d��t%0?<<6*diLI<U\i��s�����kdd}fX��������������������������vV%*]8%"?(%`q}i75idi}����c\gz��kU1?***
'86*Wv���������