Ɉb�2�-���˄VT;�rn����)�W/����|���|�k���-�`����E�Z���a;?ߖ�l
���o!($�9��Ko�d���O��V)����߳�l]���U6�J���lp����� ������?�O	\�x���v\鐋�u�Ul��َC��1��U�d�u��8d���j�@���KT:�,����p����4��Q���np�p�ӆ[<n����-���=v�n��[���� ��	���f������6�nq�l4��J�hJ�g�g3niO��+�,��L�{�kw3A���]jڶK6�d7k�-���2ꚧ0������W�}�[t6n�۸��q���-:��q�2��z>���[�:n�Ǹ����?���	�拊9���>m�h����g�[�f��#�Ym�SnMg�b�?0����>5���@�̲6w3�$�GBZ�-b�{���o����)n2����m��b��%6K�w����w��9�Ǽ�٣����̐[�>��ƞ �Hs3彡�}�=l�Ϝx�MO��=��i
�-81��5On�M�'��'捥��8��gv��Rz�,����s���eO+F��
ǩ��;��s�I%n��F��:���H{ֈ�sF<���8���d�zQ����7t�;��}��Fnp'7��[�׼�z_I�.M��M���f�y�-�3��?y��73�?;K����b�7Q���d�j�1E��D�y�4���[
#!&��0���͎����ޘ(>���3Ӂ#1k��|o���l����9HɅ�u٘x{����J�l9���l9�}�ς�*��7�0��T��/�9r������gx����S��v�o�~�~>f#o�m���D�+���l�D��y$� �	m9�I湓��)�R;
�0��Ǎ�Y� ]���*N��@�J1)P܈=�A팠�F��3�60�T鵙Y�6��/N���|{�ffi�s�/7mf��6Otz"�	���l�m<מV�X\�G}������â��{u�ޓ�n�;�F�9bA��Ḃ����Vz�Z����|��O��ީv���<�Y���5߻f���7��J��6ϓG2�������̉d)Ӹ�KL*E�T��4Lkn�bLP��N*J�)5�S�cD�FTݧb�ʖ�x�2�aጄ�����+S�Qe�9�^��Vz¨d�`_3����)�H6�K�򕃧ֵT6ye�hē��E;\�]_����J�?q��h8i^"S���+�W�Wl�b�2�2e,��Ve>]/�
��<`�jc�F��j/��y3!�e��K׍X�u������3י�^%�|!�����b���3�����W�M��ݳ��-D4h.�^	T���(���m���66#W�Ir��{��K�V�_w����
cާb���Uf�[�r�F����a*R�zG%u��*Ì�T!g�w�9v�F���1���	kc;j����r�|�[�C܎�I�s���m�ڰ45f�m�&�w��ٰ}M�T`Dי.�_Q�dg��c��7x�`��"*틸
ޛ���>�yw��А%#�-)�OY:b�eK{��S�^�M�s���@#ۼmX�z(4�a������v��R~���]�*���l���hk�}���ܧ���]._ي��C�m`��&��e�h��Ցv+�ӅleP}<(ޟ�0����	&� �n0{ײoKGl�3�.�I�<����l3KC<5�y���}Pܪ��*�֟�I��'�6%�6{�0�3���{R_�P�wMC8�����1��l⼰��L!�p{t|z^���RoT5}��ވ