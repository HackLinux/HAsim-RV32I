����^�+s���*n�p�F�>쑢5E��7���V����ׅ]z+8�����g��8	97D�!�:t�x-˛�j��iz��4ܰ��1�M���&���^x��v7ǩ�#�����xS!2w�/�$fC�r�'���/vy���y�"&��Um���p�[Rg��b�l�e���R-�4{�ȎE��bxO��ґ������UT��}_��S���«����������c,c.A�o|�f���!�ä�3Yq�����4�H6�*��܈����H�߰x�Mf���ٲ���x�5��g�"����B���ࣙ�>L=cY���"�^ԖD鎃N�%����.��F; Xj�{�@��Ė��u�^��`(�Q7���ـa[�7�f���7u%~�I%U~+s������@�J���	�k%��4ՠhk��B�X:zǬ0I��La���(?���ɨ7��o�t �c�ڴ%5ґ���&]{�Q���KF*|��Kj��0� D��=�h��/�|��<;�S�dJ��RJ[��C Ձ�)�S��Ȳ�@���Z�u���r(�WR�4Õ�7ͫ���$^��fL}���22�V91ޥ�v���,M��u���8��T>��a?H��n�B�}J݀��]w?g��e�-{M���	�esޟ%�oz�d�k����x-��V$$Q�<�����ˉ���;�9�m��Y�e�C�L���{�k�a�Y�7�2����G1���rn&gufw����Z��N! ���5��!>�]�y��"4﫱�#Ć�� ~�b�Âc�9����\6=��K\VH��-�0v�MH��F�q�k=5���݇�A:��_���X �O��:�U���i��)�N���y������)jg��ɿ�l�oH�eX��A$�����Ǖ�x�@�S���0esN�p���{�|�"�&l�3�dӺD�akH��~C�vq�����Q�f �Q;Nm�"�a/[`-�\�b�v^�1�;R�����)6I� ^a�f��t��Ai*���[��\D��� _����L� #�(�/�2�I��Mm�zA�p���7~��L�&���^�|ڑPa���C�m�N	�T�T$6H�Y���LX�$�[�%��w�X���A�!�8o7�x�
ѼYYlfql�Xl�z[2�^P��*����bsY� $��t�FK��4¯�t�K���ѯ�|������,�p1���]� e�̱ `�������<�ZE�\.(���g��]��Yi!�@E���{&^o���-"�s����9�qyC��G�	"{_u�9^n�$Y:od�XK�H�HX[m�ƙ�:��I�O0�J#SdQ2?E�ɭB���C~t�^�����%��yc�E%�X���|�>əL�T���?6��dT�������Y���'�@�Z@W���In2��E~W���;�P���hC,Xu��L��ܘ5c����*mq/]+}��(�6s?�.��][g6�e�de��"�/�H����y��^���B^ǀ�,�
��8"1�n���F�v�|�~z�����/�T'Z�*1u�m7�3b� ϊ�1	�Jx�u���$8Q�\�l�e'D�)F�b���)�]�U!�ә��D�<}�>[�LYI��(Y&�V^���t�!�i�\�^�I�M�B��Kg���^�!�;�e<x��n����xV�$�^=��A������!i^�2I��	eN�6��W���h���CX�̑�@w�kvB��B��_���u����B���/XX�|��˹8�,��rZO<#�1~�F8><����-�ױ{�L�X���g��)X�B�3 $00�Q ���,Id��h'2ޮsyEEf3'� ����6'��R��olx3Ee��,��MY '��[�&C��E�l~R0{�q���zmBU�������q��#��������aN�Q��D��t�'�_�0�b/�p-�	{�`i�}���3����.����u�� �=�E�e5��͑�8-������m�e�#���Z��|�¨�ЎM2�;����C�8#~FN�X��#(�M�E��\B�)sN�F�1�l� p��,#�u	p/��8�"����!�;U�9�0V_L
��f������ꡋ�p�}C�qy�,��Av���R���;q��e�MF�d���E0dw4�M7QR�Q�7�e��oX�4|�3n���A)�z���-��@�+�BdZN���އH'Cɝ�&��o�f�>i�����I�p�U�Kh����#%���E6������y�'�� ��G \t����C�G-v
�^��Açy��d��	� �{�y���K���S5��W��� �۟�f����\55;;�E�G/e��F�e-��0� �h����$�8hݲi� N ԟ(瀒g+?)�pC�k��������D8 ��h�@u��wO�f����ʂ��vQ�.�_
)o?�� \�}iX�P̂�j˗����"g�;XX
m����4�sJ^m0����I�Ӡ<&��TŞ�"c.�#*ސ't�-.'�4q�+��9O��.3�֪�wlMÀ=1�0��;�޴yML�o�����;�<�"�Mx������8L",HWi��4~٘�����Una���<\l"���h ։7�/����b+����x����lG"��t���VՈ�0}�e6 w����Fq&ߡ
x�S���|�\j2�F���mM(9v<��wq����������w�K��k�*��:�9��XI���P�O�d�<�x%��tE�٭�z��@CI6�"_��5@c�=�k�q������F�~3o���~�8Ä����ڝh��#���ŠUN&�I�]Ns�����6���������9�h�:*!So{�f�� ����$��ϝ�)���B�~s�O��^~�,V�-���q��&����g�,^��� �@���NV�0�u���{']?� 6i5��ҖK���Q0
#5��=<�BK�Ku8� zGA$��q*x��a������װ�c�?v���� hsO�4/�O`3��|؛�����|`�O�ȡ�=09�>1�{S���[����O9��#j�)>0@*�D������9��53(���c��f����g�yF��sN��ڽX�sg��p���"���9�u6�Ac�M�������!#9����Qh��o.��M��W
�C6�!MBS5.�(m��k�C5�w|�%�ܷ�"/�ҭI��Hx]�n�1:�ql�����뀭�%���> [y�Ey���A�H
���|k�Q$�@=�@�WWc0�*�å���+�@]�,��?L�WL�B�ڋT�<	(�{�ލ�yp�:ι% @�c#�ey�����hsQ\�أ�js�)��R��4�4�+��C���2���MɞǓzF3��;h�o�m2�W���x�@B�k�/1��@���/�����9c����k��R�u���T��`4l��x�:F+���<��@ ����U�yD��H��Ԏ�洮H����O����Տ�����%e�{j�*c�MTX#�?r��˦�MP��n�c��S��@�ڕ�+���Ñ���ߩ�*th��Z\m��6�ל��1Bބ&��.��ݺV�BU���V)��-�������pV�����2�ޓ�%'�|u �F��~u��L�>v�,��^w�r�V��������+`b������Whd%M�`,1�'BհvB�AZn ���xk�9����?����e_h��&�"m+�E� �04�˴����F]|��~���g�s�п�Q�:�v�=��?9 �h<���>۟��&�8��9�]��sZ%�Θjm��$���p��!��jmƵ2������i,ݪl��Gn�X�V)���V	7YТ��w��t�����ĹMe;��ɣɈ�-8��X���fq��q�����䉂��ƽ5-<"� #nn~�j��˄���U@2��P�7� bD��$�8�uM>��9�19�Z�;fZ��O��e-��m�ڹy��=�Q�(���4{K����)Yz9'�;G����=����[m��,�Go��/B^����Q-���_HW�Т9E��ϩ�����n�M�e^�8�}B�t��צ�<��ӹ^�uBf�)���ѷ�AI�^���*�K8�z�gavQ@g3T"��k�@ĵJ��7�����N�P�ȕa+חQ��q��xkc���0���� q\�~�z��|	�������`I��<l�'���ؒ�B��tq	!~���Z*-�G)߳�m*s �_���r_���p����	��C���X,�3p�u�]~��<�"z>Mw�3b	߆�bߚP4�Ѧ�U�3��"M+���;�e����F�1�}�ظ���
Y�@���T�9?	���+:9�z�;��+{1�F�f� �|���>�/Z���9W�Ck�;�MND���/����amEݡ���،rAU��K�t2��ѳB�lcƭqs�f����s��Ȩ<1?N�Z�C�~�]Ӹ�i�)9�=9��<ء�!�����-)�^��×ﴪ�
�^F4����,$vO�&����S�0?rj#�0Q�GR��[H�b�X�Q�G����M�\)�	�f�רv�%�`h��Ӣ�<׉���Ea��p3'�?a���UҘ�����*#�y?�ZFr�5�5�z��ىy�_�J oz.�
/�)�dږ�F:���a���=8��4��r��
�{I$]L����R���%n�GlU�����a��[J,d�4��t�i�����{�t�������9b��uCA �Z��31�2�WS��u��O����8t7�x&H��I��8�z�ս�6�Xn���X~�W���F<^K��׸}\��>�VM4�(~���tP��K\EX�e>jq��-h�<���V¬��b�ˮ���y��T������F�5��|�{NrT����FH����5�2ؿ�1�B�d?�`ܘ ]�M4[oh���u`��N�1��%���A�L�g1�C���\����H�<Q�g���0�bA��	�<6�9�K���'�=t���Z���*�@l&�ޜA��u Θ�_��8��uW�?��{8Ū}ش�8�D���Q$����4��q#����T���h~%����������6���[S����~!\BP�?!h;R����d禆U�I�'b�w��;`�1l���݂4;swU~����<V����7B8��:"h�!o~I�/�	%�n��tw��V�Y�O2�j��|ڃ���iT�S�VӬXh���0�pCz�e��{�C� d���`ud�a�c�<�Ŕc�i��t�)�;��6��8�<6��˦��`D�ptf��ǔ������/e�l/;J��1���N���h��΍G¦�w0ŝ&m1��Ah'���
̡׷H�|tZ"�'^+wRF�x�<?v�H�GHA
�p�X,�X�0���Ņ?�_��fe������QƱ��犩)��B�h�/�o��R4E�����8EG_�3RxA+�ԝ�j�znU�Oo�5���f#l_��[���q���\����Ҙ_��������_	�_��|Gugޞ�b���b���b/Oh�ghqToh�Twh�UhqVh�V'hqW?�]�cm�-m����`�? �T����mgP=����T~C+��Y��Oj978��K��g��j����ސz鷿3�D���j�Q�a5��ߨ�`�_T}Pןu���
|���I}�w+��~���̪��8�J���m�*�ka�Q����T�io0���F�U=MV������n�WW�x�f����
��n`C罓W?�?�]�-ܥ�ݞ¾z�����/�����;����Qu�D�������<����; �@KR_c!b��!�uC�ƏW�6*�qj߭���L! ��a�����Џ!ν��c����o�����~����P,��ݘF�������ER���R�X���d��;�d��y�ɓ.M��b�O0�}����|��C��ؘc��Z1�[�QY���0l_��y6����E�m��uu-��b�j���p<���S���a��_���=�[��L ~0T�~����c���G���XK+�\kh��o�E�d��݋�%l!����a����A_r��̊�L8��_�q�:ɗB�W��(I:���b+YPC��*Wӓ\��|T�p'�/�z���3aP�Q�8$�IQ_�����u��N&��DXxuk>g4XHs���]]��h�r��3[۴9�6�<��/۱U�0n��i�H4,�P#DR��۶�3;΄:��N��^�GO��uw&��k��(���J�o���Y�+Gqy�=� ��a��_<��5�F�T�(Ep��1qjj/���c�{;]��p:syp)D+��H�sN�1қ��W�������v��c_�%S��j逋0�S����P�`%��E
���E�b����C��'3�+�h�)�ƺ�`�[ނ͕(ޒ�!���h���X��=�Tݛ��l��ˀ&�5D
�a������Y��o���刍}�j�3K̀1U$y#����<��u@e�A\�9o[�e-54�V5 ��H��ޛ}����3Mň�L���E��~����;�����C$x5H%��f����K�``��(-G�w!��L8S�D,c��Z8C6K3q�pO0K8
���M~N0�l��r�s�P+�j������Z!�A�����d��I(�KU�M!�ͳ� ��TA9T�L��Z	m�S%Jެ`�W׉}��3�ɞ�|��=�"h8Pi݀�c�
���v���;q
<�g���b-��N�o�s�6�@ƾ⁧��6�w�t$���N�D�N�����xF��T`�'�}�?#S�65�4�p�1���qqp[��*ߩ�P��{-��l3g_��hB�������Θ<��D������l��$'ܨ�4!��пNo���Z�>Ǩ�B���m����!���o���?��_f��~3ӎ���FR �㌍�.�ʲ�Yf3V�OA��5�ސ��j]���H}�Ү�1A~?џ�±�i��!O�Y|-˽�<�>���<J"� 
���\��څ�t�yq'.�7^\��ƥB���ς��^{z�ʱ���؊�t�tc�C�-��d�n�g��S;��<լ��i�:�M^^ؘKf%��.tI�"y$Ĳ�f�Q7Fp*�9��/�O :�v�=�T���*kLR�&dC�aLH��4|_����K�呆A^L���94�@���q��KdO8�{Li.u��\(J�u)m��)��H<���iy�+ i}p�H��ʂ���N0/� ��Ag�m��D �&Yᣪ��V)ʖ$����v!��*�IQ�O*���$��L�x�K#�����m��<&����f�&۹J6����y��kC�M���o���`��Pưm�������[��Xz-�G��r�V�gh܉Y$G�k�b���x�s���N�'���0�I�	h_<ů�af؏�P)�Gآ;��EO
��en���O�t0WG��y��K�	����X���u�5����]�����J�`5�/�;�<"4G7�gjͪ����h�%M���M���]����uQE�#��#�^tf�Zo�����S�O86y��'�<f��4a�(���ލߠ��g|�=�T|+jz�`^��8M�t��d��gY*]�1�o����*r[]Z��K��)M|$p��n���Mel'��k�mIV�uEr��牞���H-�Z�)C������D��E	F'��:��@Q��7��2v��RF���N�r)������%>�ӂ��;>������R��7Ur>y͋�5ᐊ���ky�ݢƤ�Ƽ^�t�Yj���g�jr݁�\�����@�1�c܉0KA�R ��-����(�� ��^)5&#,�W���;�zv��Ჾ�Ay�e��H������`�;��V�)� 9t��]���A?�������)�y��*ރ�I���$��td2�RY� .CelQ9����|�-"t{�|�/��Xj��v
�i��&d�M\�)c��S���������s��E1�OcT�È��ȭ=V���rBJtԂ���T`�j�h}�bǺ���v�XL&���q#� ��B�s����]��az���v�)��M�Qb��uhe�r`���1���K	ʪ??�So`�a�z�HS�+a e5*a�j�n�G}�t��T%��P��hZ�em�O<��H<����]�����S¨���B�5C1������o@��вzK������uo�;����NH�^���~b�	�w�e@��5�$�z�і�X��B@����}�O��3��6U�_�*�#����f�1�?Z=tS�?���lNO���o<n�w�.3z�U�G9�=��ץ�\Q��{���m�/�8�_��(&@̝��q�'7�h��*��̓��>	��5�.&��ѭ�/,��������v���-�@�9��f qy_`
5
��L�ƿ���w=G���߱.���M��K�NB�5Qť��QcX�Rj	N�����O8�X�O���-�?��	?�P(��p<��z���	�ɱ��`�B���'G�2��#J����=��n8�W������$*�"��6K@���/��%��0+_=�k��R������q�UR��~��;^�|�De��O/�z�&>����}�GT�nc�F�XBAJG�\�O���P]k5/�Z�Ѧ����ʨN�6S��;��vP��Nd8�e�"���$�͏q�v�x�Uh|so�)�x��,�`?�Q�Lѕ�]qfQ��'��B��=�G߷d��%�u�Q���=V�i
ﶡ�xT�t��'�J'#�S۰��~z<�Ň�U��6DR"|���[y�T�0���԰�v�U��"���x�3�O��r���{�S�#�؉�m�ŉ�o���5�"�Cv ��@+Jɋ���֢CM�i7ħ}��P0Z��3ȭ���=8`�I/���@G�~��K鱧�B�T^�?/��H ;��h��u��o�ƷH���KK2�r��61���P����a�?|X̶w�cH�F����p����1�����hJf"������a��XK��cdv�R$lNٱ�('Q���T����W�74��[+O�{�W-�^IX��KT���~E�j��<J��7l
�d C�1�a�U�x|c��&kې���)~d���>l-�e�C�A�SZI�|�ou(�c;�c7�x��g�v'�s!^��}B
���@;Ͷ_缾:YO�U����<{Fm�4���gǻ�=�8�&�wq2�[o�2/��۱��b��5~b�
��N������3��֠��������1ր̚Ж��j@���r��8Z�c���c*�ݙ����f/!$G�q�1���DN�m]��+/!��a.�V��/�Lݧ��������&?�y~�56�lyD� R��V���x���@|�f����m�eykˌ�E�u���*L�Ɗ9�ҝ@� K����ݲE���(R��#puؑ)�2�p�/�W^�pFJצ.|�\W�^��ko#tPz�	����