import Vector::*;

// ******* Project Imports *******

`include "asim/provides/hasim_common.bsh"
`include "asim/provides/soft_connections.bsh"

// ******* Timing Model Imports *******

`include "asim/provides/memory_base_types.bsh"

module [HASIM_MODULE] mkMemory();

endmodule
