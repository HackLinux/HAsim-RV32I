��������������uu��  ��22��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������@@��  ��[[��22��  ��uu��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������  ��  ��

��

������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������  ��  ��22������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������@@��  ��  ��uu������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ����    �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ���    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ��� ���    �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���� ��� ��� ��� ��� ���    �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ���� ��� ��� ���         TRUEVISION-XFILE.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     