-, 0,*�/,+/--.,,,*+%#$$"#!!  � � � � 1F.?*:'8,=�+<.?+<):*7.5P�?Le$>Kd9Fc?OmEVsI^wKc}CTs;Fe2<Z+5Q07R1:S,2F-8Q/:W1>];Me@Sd6DZ=d{=c�?e�Ep�?d�9Zs4Tb@bnDhtAjwEl{Bl�=f�;ay5Wo7Yu;\{6\v�:_|6Yv5Vm9^q:br3Qi%.K/8S/:U7He6Ff2Bd8Jn/?c8Jj3Be/=_/>.>+;'83DK6HN�7IQ}9LS;OW>R\>RZDXbPhr\w�v��������������&9V&8R*<T&6T%5U'7U%7K*9!/I':]%7Y&;V%8K#2G(:P*?R'9M*<T-B[/B]*?X'>]&B\%>U*AX8OnHg�No�Vx�Wq�\t�f~�u����������|�����~��g��u����������nzzouwRbdHffWwvc��i��`|�KawN_vWe}[w����~��}��q��`u�j������³�����������������������������������������������������������qy�y��m{�t}�py�v~�al�is�v�����������bd�bf�W\�HDjSJnRJjZQs1Oa4Vh>cv?i?h<f~<cz:]t<b|?j�@i�� � � � � � � � � � � � &$%%#$�&$%&$$&$%)'',*+.,-0..1.-�.,,/,+.-,...---,*+/-.+)+�*(),*+,**,*+.,,.-,-*),**.,,,*+.,,0-,,+*,**�+*),**+)**()%##$""!  � � � � 2?.?+<�*:Q*<,<-=1D,=,;$+D3@Y@OjBOh?Le?PkEUoJ[tGYsDWz?Lm9C_1=W1;U;Ha7BW*2H*3P1<[:MfAUi9H]/<U>j�>g�<f�Gt�Dn�>b|7[m9Zi<^j@epIp@h�;a8[v6Zt9[u<\x6_v<c~<a~8Zv6[l5]m5Zm&A*4P.;T6Gb4Db1A_:Or4Eh4Fh6Hl4El+5.:1=2B,:3DK6IP7JQ7IO6JP9MU;OW>RZKbk_y�u������������?���'8U#2M .N%4W%5S+J"1H&5N$7V&;X$6P"5L&8H*<N+>Q)<K&6L0Gf/E]*C\+C[+D['@S';K-E[;[kBgxHk�Sw�Zy~ax�r��v��o�����|��������u��z�����������_ioSekWek9RY?]eSmwx��j��as�`u�h��Zp�h����r��k�cq�h|�j���������������������������������������� �������!������������������z��~�����ik�jp�Xb�Sb�OW�nu�w��������Z[�RT�A=ePJn]WwWOoa[}@fx@l�?h;f}<dx;as=d{?i?eu� � � � � � � � � � � � &$$%##&$%�&$$'%&*((�,**/.-0-,�,**�,*+�+)+.,-+)*�*() ,*+�+)*,**/--/,+�.,,,*+.,,1.-.,,+))�*)( +))�*()$$$" !! !� � � � /;1@,<%5(6+;-B�,=40B2@-7Q)4O4@\CSmBPj?LgBRlGVqAPi?Lk@Sv;Ig5@]0;T5@[ARk/:S (D)2S5Fe;Qi5D[/:U%0MBs�>m�:`~;i6^n6Xj=^s6Wl4Uf8[lInDf~;Zu4Nf8Yn<^z<`�6Zx:_|?fAi}8Yn3Ti8&/L/;W5E]�1A_6Il6Ip3Gg4Eh9Mu-?,>,;-:0>*72DL6HP7IQ8HN7IO:NT;OW<OVNdjk��������������������&8V"2P$4T$3T)9U�&7Vj&8X(<\)=[$5N0E+?W)>S.DX%6K,>Z1Da/E].G^.E^.F^*CZ+HW2O^BejDjiJuxIlo[co������ew{dy~v��������}��v��������������Z^`[wlY`i7H[;Ja]w�e~�k��z��z��f��[p�i����s�lpvZctb{�i�����������������������������������������������������������������������������:_p���������ac�KR�EU�GS�SY�Zd�fo�s}�el�W[�IKwVTvfb�c[{b\|dd�An�?j�<ex?iy@h�?g�<c�� � � � � � � � � � � � �� ���� � � � F!'E+:,;+:)6$1(4,<.D*=+<8E`1:U,4P*4P4A\DVrAQk?LkBRlCQi9F_;Kk>Rr:Ff2=Z1;W6Cb0>`#H#C,8Z7Ii2B\+7S".H)H=j�;c}8^x;f}:br:`r=ey6Yp5Zo9^u?_w;]s6Uj4Mb;[o?b<`�6Ux8\x=c}@f�:az"9"*F.<Z4B\1>[2A\0@`2Dh1Dg3Ee8Lt,=�,?+<,:/;+62DL4FN6GP8JP:LT;OU;NU;OURhlw��������������������#4M-L$3V)9Y/A]+=[*<Z%6U$3N(8R%6O%7S)>S,A\.C`+?],B`,?Z+@[/G_4Nd,CX+FY%IK>\d?\aAihCbgTmz~�����|��j��l��������y��u��������������}��brq[igL\bN_hWo�h��z��o��w��~��q��t�����q��hqth~|jw�k��U����������������������������������������������������������������������µ�����:_t?_w���������jl�PU�:=|AM�HN�PU�KOyEGqX_�[`�QS}WZ}fd�f`�e^�if�os�6\l?h?e�=d�;a�� � � � � � � � � � � � �� ��� � � � �-;V.>)9'5'4$1+9.>/D)<9Hc3=Y/7S-5Q&.L0?^CVs?Ok;KiBPj?Me4Cb9Lk?Oq8Ed7C_3>]1=]"L>$A/;]5Fe,8X#-M(I'J6_v8]r<`t?j�?k=g{;ey;au<bz=c{7So4Tl2Of4Nd>_v?d�:_�3Pq9[w?d�Bi�"*B"*F0@^3A[.=X2AZ)5S+9Y/?a0?b8Mt-=/D0D1F0C0=1:5A2FL5GO7IQ:KR;MU<PV>RX>PXSgky���������@��������� 4F.J!/O&8V(9V"3P$7Z"2P&4L"0D$4J':U,A\/Gg1Gi0Hh-C_-?U/G_4N^/Ja-I[&DL/NS7NY7LW;QeOe}j��������x��fzut��������������������������imuXgrNbh?UcPhzl��y��q��z��t��j�����}��g��h��\qz^nxw��d{�Usw�������������������������������������������������������������������<bz6Sn3Qi2Of������mn�VX�<<n64fFGxV[�IJq96\KKuah�SUMMqRNp_W{g]�kg�su�=f�<c�;a<a�� � � � � � � � � � � � ����� � � � .:/:3?0@*9%5"6$7+?0F-C:Jh3>]/:W/8S,7P'J1>[ASs:Lj5Ee=Mg:Jf6Gd?Om?Oo;Je?Le;Je-8Y><%(I0>^4Cb)4S%3U'L$0T4Yl8^lDlvFq�Bp�>i�:apAk}Cl�Ad}9Tk3Li3Lm2Np=b�<c�6[~0Mf9]{Ah�&0J%-I-;[1@[,:V7H_$-J#,G,<\/?_6Lt.:1D2G3E6K6G7B7>+9Y4FJ5IO7IO7KQ:LR<OT?RW=PUPdhs��������������������!/=+:O*:T'7S%9M"5P#6Y%5S)9Q%2?"3F$9X/Gk-Fk*Ef'?_-C_1G_5Ma0HX,EZ1L]3NY5Ma>Rf8Kb:QtWv����t�����bz�m{{p��w��|�����������������r~~Z[hRdvPbjHYl^{�w��r��r��z��x��{��y��~��w��j��`z�ats��]p�ey�����1����������������������������������¿��������������������������µ�����?by7Ri3Ki3Lm4Pr=c����v{�WW}==i/*T;8`TU~]a�PPxTT~bd�_d�IHn:2VLDhbZ~jf�qt�~��<b|<d�� � � � � � � � � � � � ���� � � � � ,=*6-91@,=+:'4#4(;)?+C,9X2?^,7V,8X0;V*6P#'C3=Y?Ro5Hg4Dd:Jf�>Nh<?Pk<LhCSkG[s=Lg*7T;#E'+M1=].:Z+9[(7\"2Z+8];`s?ewClBn�=f�:`z8[l@fz?h9]w6Xn3Og2Kj5Qw7W9X:Y|?`uBh�*8N'0I+8W/<W+7S9Lc&/L#;)6U/>_4Gn/;0>4D3E5H<U!>W$?T-?i2Bd3CI5GO7KQ9KS:NT=OS�>PT\FX`Wkqg}�|��������������'1=1BW/A]&3R)>S#;[&:X*=X(:P5> ,@(=\-Gk(Bj*Ad(>\,CZ/DY2F\/DW5Pa:SfAYoDazA`�Ib]��n��~��u��h��\|yewyh�s��r�����������������bw|N`lVk�f��a~�o��o��q��w��t��{�����������p��h��WwwT_lu��v��y����������������������������������������������İ���������������������������8^v6Wl2Mf3Nm5Qw8V�9X:Zzt|�WX}FFr;7c9IGifg�jl�or�ed�kn�WX�A:^E@db[�gd�op�z������ � � � � � � � � � � � ������ � � � � 0D.C)<'6)5*5)4)5(3%2):*1J#-K+7S(1P*5T/8U/;S*2J(*F2@`;Li1@a5EeAQkCTi@Qf?NeASmK`yASo;Ke.:V&F#)K'.S-8W#,M*:^'7[.Bj3Ei>ax?e?h�?g�;_�7Xw6Wl7[m8Yl7Xi9Yi2Rd2Nf6Ut:Zz;]?`�Ll�*5N)3I)4Q/:U,8R>Qh'/M!)E'4Q.=`0Bf,:/>4@4D6J;O!?Y#AY.@l6Hj+8W2BH4FN6IP7JQ9LS:NV;NU;MU=OUCW_H]fax~�����������%.?-B_2E\.A^&=\&<\(?V%:K&;L!3=$0F+Ba+Ek'Bg,A\'?U3J_2H\2I\0G\6Od9HY9GU5Ia>`xNr�`��x��u��k��Se�}^vxNk|_�����������|��}��������i��[t�^{�s��k��i��m��k��o��}��{�����}��s��i��cuft�fx�i��}��}�����������������������������������������������������������������������������7Xi9Yi3Pc2Oh6Ut:\|;]?a�Ll�z~�QSsMOwGFt74Z?=[on�yv�||�uv�np�ou�VV~TS{ab�kc�hk�w~�� � � � � � � � � � � �  ���� � � � � W+?.C+?(;&5$0$,(,(1*2)3*2J&.J(0L)3O+6S08T,5R-7O,4L(1T/>]0<^2Ad<NnCTmBTj>QhARoEWq?Pm6Fd;Ke/=Y"(L$+P-7W&,J&1T)8Y,=d@U�:Mp=_{<`~=b�=b�9Z5Su4Ph-K[1NW7U[;Ua6Ud4Vf7[m;au>h�Bk�(1L(0L&0L-8Q0=V=Qg)2Q%/K&2R.<`,:\+:,:0@8F7I8M!?W!>W2>d6Hl5Ba 72BH3DK5GO7JQ:MT�;OWz<OV<NV?S[AV_Tlvk�����������)<U);U*=Z&<\#8[(=\*?R&8B&;H"7D-?[1Ii';e$;Z*=X2H^8N`4HZ5La3GY3DS0=J.8D/BYGh�Pt�c��z��b��w��w��\ivm��v��������y��i��w��������q��k��x����t��g~�Uy�s��y����������}��q��t��x�������������������������������������������������������ż�������ŵ��������������������������9V];Ua5Uc4Wf7[m=cw?g�Bi�Om�Cm�?i�YTvEA_PU�ZZ�WW{ml�~~�}y�~|�uu�kn�gk�^`�ad�d`�hb�� � � � � � � � � � � �  ������� � � �  &8�+<V*;'8'4%-%*-5)0*4*0F(.H*0N+5M+5O2=Z/8U*2N-5M,4P'1Q)4Q1=_:Il@TtATo@Sj@Rp?Rq<Jh6Db8Hd:Lf1<[&-R.6V6?X.7X0?f,;b6JvG^�;Ko9Yu6Yv9^{8]|5Yw4Vp3Te/MU3V];^g6PZ9bq:jz8gt2Zj:dz'1M(0L'2M,5P3AY;Me(2R*4T$/P,8Z)2U'4'6'81A%CO#@U!?W"@X3?e2Cj:Ij'2M"'D2BH5GO9MS:NV;OW<QZ�>RZw<QZKbm]z�s��������'5M':S&9T'<[&8V,C\,?P,?L"8H(<P.C^)?_&<`&>b,Db3H]2GV.CP,>P3CQ,6F(4>)9?'<[F_�Wy�c��f��t��q��m��cp{m��~�����y��l��\x�t��������l��x�����z��b��PgxNg�m��r��x��~��~��~��w�����~��������u�����k������������ï�������������������������ſ�Ļ����³��������������������������;\g5OY8dt9l{6ht2Zj;e{?i�:Zr8_v8^n6[d8^jB6POMmY\����kh�sp�|y�x�db�^b�`i�fk�]_�\[�� � � � � � � � � � � � ������ � � � E.9V)6):*>)<):*6(2)0.44>#&;(.B*1F+1M*2N(0H/:S4@\,6R,4P.5L*2N%.I+5W7De>QpCXw@Un?Pm;Oo9Jg5Aa3A_;Lk9Ii1=_+5W09X6=b6Dl9Iq1Bq<P~K^�9Iq6Xp7Xw9[}6Wx7Zs9Yk6Sb6Yb:ep<iz5Vg7cs:lz9hw6`p+5Q'1M)6O,4P5C[9Ja'2S,7X$-P�+6W%.'0'4)80@!>M$CX$E^2@h6Jt:Lr1?_*2N&+B3DK7IQ:NV=QY>SZ?U]?V]?U]�?S[T>RZDXbLclTqzo�����&4N+9Q)5G(8L)>Q,@X,AV)@]*@X,=P+=Y'@a)Be*Cd2Jd5K]/IS-AM2?L'1?$,8#29#0=3JcLk�\~�e��r��s��e{yb�~o�^{�[z�~��f��f�i��r�����s��q��s��s��f��Z{|Ylyh��t��e��m��~��w�����������������~��������i���������ù�ǯ�������������������������Ŀ����ñ��������� ������������������<ix3Te9eu9l{9fw6^n?kBm�;a6\t5[m6[j9Zk3Pc^Sw^YuZY}fg�kn�aY�pm�mf�^W�DD|SY�gl�be�� � � � � � � � � � � � ��� � �� � � � Y+<)8+:,=)?(>*<)5)1.76?*1D*0@+2E.8L+2M'1K/:S9Ia0;X+4O-6O+4M&.J#+M-8Y;KiAWwF\|ASo<Lj6Hd+6S,8X<Nn@Ux=Mm8Ed*5X-7[9Bk>Nx@S~9IAT�I\9Ju9_w;]}:Y�8X|:[t;Yi;WaAhs@r�>p�5Zm7`m:ft;j}/<U'1M+6O+5O3@Y7H_&1T,8\$-P)4Q,8X#1%.(0(3)60>6D"AV6Jt=U�>Sz:Lp.:T-6O,4H6GP:LT;OW�>RX >RZ�>T\X>SZ>RZ<QZ=QY<NV>RZUqyk��&6H)3?".8-8&9J*?R(AT'Aa*>T*5@%8U&Bh&Af/Ha1Ka2L\)=E)9A*6>$4:07/<(6J;SkMg�[y�e��m{qyxcss^�{\nv\o�l��u��g��_v�w��{��w��i��p��k��m��^�}S^kn��s��r��t��v��z��������������������r��z�����w������������������������������������������þ�ſ�������������������������Ic�[y�7am:gv;h}:brAkDp�?h�8^v8Zn:[p5Qe1J]1H]4Phwy�li�MNu[_�ZV�WQ}RNtWNzA<pDCsSY�qt�� � � � � � � � � � � �  � �� � � � � -;.?0>2C0E*?,C*?'7+229.8L.5J).?,5F/6K*2J,4P<Pf3A]'1M�+3OB$*F!$E#*M,:ZAUsH`�H_|?Qm7Gc!)E%A:NpE\E[yBTr<Np&2X1>g>LxFX�GZ�?Q�CV�J\�>Q|Cl�?d�8Y�;]�9Z{:Yl@_dNt~Jv�>k|4Zf6Zb<cn2A\'1K'2K+3O0;V5Ga%1U.<^&1R(3P.;X!,$2&2(5(7)8/>3A;R}<R~CW�>Pv/;]2:V)1G1:U9MU<QZ�?S[~@T\AX_@Y`@W`=T]=S]>T\>RZ>QX>RZF_hPjr&3@%/5 3617#2C.EV)A_'>e+@Q$-:#8U#<a,Ed.G^.FX+CS*@H+;E(4>$4:29*;1H_E_uTq�_��m��r�zu�|ey{cw[r{`}�t��w��g��v��}��t��e��n��u��m��r��n��l|�`~�i��}�����������������u��z��������z��{����������������������������������������������������ĺ¿�����Ŀ�ĺ�¹��������������>NlSk�_w�;dq=k�8]tAj}Ep�@h�?d{?_q?Wk0DT2M^7Qc9Oa<Uj<[ntu�]\�EHsW[OKw@<hD<fGAi93_DEr� � � � � � � � � � � � �� � � � � L+7*6):/?/C-C+@+>'8&2(0F2<P/9O-3G',A+1I.3J*/J1:W4D^*5R(0L+5M"'B;$(J!)I1>[IaIa�C\{:Jh*2N1+6WE_�Ib�JazMe�AU/<g:ItEV�N`�J_�AX�FX�M_�>Oz>c�;`�9Y�7Yy4Tl4Td9]gAekAgo>bn2R`6SZ5E](0H$*B)2K.7T3E_%1U/=a&2R'2Q.=X#1'".&3&6�):1D=U�=Q{E\�AR},8`2=^&0H4=X19U;NU=QY>RZ?T[AX_CZcD\fBYb@W`?S[>RZ@T\CV]BV^�@T\@+;C",4.2#3=.CT2H^)@_%?]&;J!.;0M'=_/C_0H^-CQ(>P0BL->E!+3!.9.<(7L6PfH]rWr�a��m��htp_kkMYiLcj[m}o��|�����x��|��v��{��z��r��^v�h��u��i{�Tn�Oq�g��r��������j|���������~�����������|��x��t�������ķ������/�����������������������������ɴ�����������������������������)2ECSqM_�Vd�qz�6]tBj|Eo�=g�:`t8Yh5Ra2O\7Ri6Nf,BR2Rd6Wn:\t;a{ji�OPyIJqRW|D<jC8bD<`:6\� � � � � � � � � � � � � �� � � � 	 4+".&3&6'8):'8&5):�'8,>.C.?-9*4.7+5'3/;.;,=-C(<%6&-H0:R09R07N+2G$*F�*0H+1O0=\-:W,4P,4L#+C7&+H*4P (D5B]E[{C[{;Mo2;Z$&D;7EiKb�Of�Vm�To�DY�;JuFW�Nb�Qh�Ia�DY�JZ�H\�6Hl;ay:_~:[�6St3Pg2Sf7]o9]i;`k;`o2J\-;Q'/G 8(1J+3O4Db&2T.<`'4Q'2S-:W)<$<0!0%4'8):+<=U�<Q|E\�BU|'3a0:^%-I09T*2R(.H:NV=QY>RZ=QY>RZ>U^AXaAWaAW_?S[?Q[@T\@R\?Q[>PZ?Q[#4=$,+6,?P1I_0F^'>W#;K$:D$:@%8S,?\/E]*?P-@O,=N-@Q%9A'5 )<%6K1G_?YkKaw]�f��o�ageOOQHOb_jhz�x����������������y��p��%p��RgvZv�`t�dz�Tj~a��x��y��x��h{~[`mx��������������z�����r��i��^p������������������������������������������ȿ�ū������"���������������������((0F<HhCS}Q]�\e�ow�Dl|>f�:`z6Xn4Vh:]v<]�:T|0Kf3Oi7Wo9\w;_{<b|vx�aa�FFnMPuHGoC5]ODf� � � � � � � � � � � � ���� � � � � � \$>"7"1$4&6'5*7)6$4):);)</C,?*:*5-5.8-7$-,4/7-:/C(<'0M&.J*2N'/K,2H'-G$+F'/G(0L/;Y0@^/:U-6O-8M$*B(.F-6Q$,L#=,7RAVy?Tw/?_.5T" @+1SCW{Of�Xq�^y�To�I^�L^�Sf�Um�Nh�F_�FX�G[�=Pw-9e9`m9_w:^�6Pv4Pl5Wm:cz4Yn5_q8ar&0H(2H4(/H)3O-<[&2T-;_(4P'2S.9V,C,G(F$>$6&5�'8;Q=S�BZ�CX{2Cn+4Y'/Q'/M$+N!%G'-A:NV�>RZ	=QY;OW>U\AW_BX`BV`@RZ>PX>PZ>RZ�?Q[=#7C+7$4D2F\1F[)>U#;M&=J/DO)<G+CY+@W+?S,AR/FY/DU(;F!2? .@(<H6IZ;Qg:StPk�Yx�\�e��^vjVdb_tyk�����������}��������s��y��}��e�|[fwMh�QbwZgt\izp�����z��~��_pw[jwv�����������������x��`��]q�c����������/�����������������������������Ƨ�����������������������������'!5,7P8HhM[�Xf�O\�Zc�]b�;[8[|7\yAf�@c�>\�9V�:Rr:Vr8\x8[v>cx<^t6Rljq�`c�JNvGIsE;e� � � � � � � � � � � � ��� � � � � � (A&="1$3&5#0�'1%1)6+>+?0C&8%1'1.:.>,:$/*6,9,<-?-5U'/M�!(G;#)G'-C'-A'-C(.F+4O0@^2D^/:U-8Q,8P+4M*4N%/O &D-+2QKa�<Or7Gk.4T/8]>MnJ\�Ul�]w�i��To�Sg�Sf�Tl�Sk�Ib�?U�DX�@S~&2`-<m:^r8^x6]~9Z6Xt6Zn7_o6_t8^t&;(1J!$=&-H&/J&0N&2R+9]&2N&1N-6U'<*C�*G)E%7$4&83Gs=V�@V�F]�;Ru-6['2W(1R$J $H,4P&*B9MU=QY<QZ=QY>RX?S[@U\@T\@SZ?QW=OU�>PXE>RZ?S[>PZ&8D%7E/FW)AO+>Q1I_)@S,CX/DU*AT-Ga'@S'<M,EV-Da.EX&8D&9L)?U-DO5HY?ToFb|Rt�_��b��c��e�{hrtl��i��~��u��}��y��u��t��m��u��t��h��Vmxa{�_u�dz�i�������f��{��[kq_u����z��{��������~��aouMai\jzk}��������������������-�����������������������Ʀ��������