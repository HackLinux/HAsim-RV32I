��&/b�G��-�$��Ep�A��+��c���l�i���9GJ哠IRnG��#S*-{�X�;#iQ�i�X(�-��w�,H!���G����5J0�������db�T�n
�ד:�����'�_���3�� ⒅�ݹ T������D	}s�u�F��֪�Z�T�fxX_�(9�T�" nmL�� <Ū�G���)J���p���6̮n�Q�A^�cf�Z]	>��s���ja�����%�/�>g{\!�9m��KJ�G�Hp�8�K���&�b75�l6?�J���F�RML���z�Z�-x�����]~�6,�d{>bN�W
E�Ѕ�dOZHS+�-���_�7�vS�U�4���]n��O�{a0.���L��\�Ķ|a`�V�>\Y�L�2�O��Sp�M�PpǛ\�n�Q�Y��s�c��n|'4cO�T��C�0��ݔ,���قbO&��Y�&�=�j���㯧�W��ɟ73-0q��WG�����'��0��@Q
h��������Vǉ����S��7r��|�N*�v��$����'(S[tZ�F"ws��'E�<�Ϩ�x����O�+P��c��{���kֿz0-�m���fF�����*�1������e6"�}nbg��"KnB��� r&`»*��VpnUUA�F5k$L�7?4Q��"�H�kH�ؒ�w�U�{&{U��87�Y�:����G�E=�c�Q �Ope�C\\��H.�</��&Q=�e��"��g�'1���d]��Г!��C@7��?����X��Ĉ��b8�a��a	 ��Ai�O���8�%(� �r|�QV��
���45�J�� 6|��2v��4V��x��e�f &�}}��|G���X��Ƈ��m-=����]<�~b�%�Yܦ':��$�T��c�T��G�*��O7�7�i��ύ��f����� P<;�mW $V��	��*Q�7~o$F��z�k����޴DU&B!US{QH���:�
��W��B"�+Rt�*�_HE*֓��I�Nb�F��)��!)�t�gAUe����]��po9�?h,ί�9���`@k��Ɛ���dЈi"� 2�����΀�1$₨H7@C�U����dnH�X;]b|�\��g<��4�8r�l�)��6t�*�s���q��d��`�6�>���/@��ѯ��A�w�Y��2�Sy!�e�pȈ�#��pZ2�5��95V�-�W�j7��/�C�8�t�}�]��L�87�����},! �ɂ�H�CՏ�a0G"�'���#l�B�J�����褲��V��AuB���:o�.j���lj���u�	���.x*+u����*_F������r/�Z��臯��i��E�N$M�!?L�­9�y���S֮��(�����	T�,@�Js�N�{�k��+������R�d����t�ےkXw�k��x|��1P������N�I��B(?��^5j�C��WZ,\�c@!-	`8w�`��?�$��V��n�Z�_{mQ����a��]=����5��Ӎ�q~v2��4pĦ�hD8K��z�)�W�wIџ��&$��x}	{Ϣf �Z�DJ\P: ����[܇A�^�]S%�f*��[3�O����,�^�=(w8�9�I.��-����,�H�-�Ζ�#\��|��6����9�wӶCy!v��r.F��LMN������uC�q|��G����2�T��=;�ڳ:��E�+2�ttMNQ
��<@+�p��,7Ǐ��kLqTW����B�X��j���!̐�M������&���ؿs�}|H�IN5��x#.�;��ƞ1)��r��K�����*d�x����D�<it����U/ۯ��t%$\ñ��1����X�eaq�B�,G�*�"��s���H�߹b	��jFN�U�j0���W�e���]Xbƛ�J��b1�m�b��S�>tRN'�U��w3�Tv�xW�<,C�XN9�C^l6������?�7(!Ņ+Lg��1�\?c��@p\�'  �և�{d:,��Sb|�tS��!��c�^. �v1b��fE���B��z�Uك���!����d�����Q2L�ا4g���#ٴ�/�'y��s��l��G/Q5ԛ|�.Y�N�1�17�7,���`j`�,����Ĭ��x��0*e䕄�����hp�U�k'1��.���k"���h�Q�3����k1f^����$��C%0�?�X�í1���l`47��V)J�G+�B��/n��.�q� h�r�T���N`	rq��'�P�u d��O�����6��}�lQ�!������u�ǝ.<ձ���=�L6�b�+[y�zO5���FI)��6�-�)@���3��.h�t�/�� D�;�ō{�}ܙAUQ�"��H���a��\�w�9qw��g[-�o߻�~v����f���r�.~��ɞ�,B�U���]���O<��Ο��S�xԎ��'�r���;O��&fw��ApR;B6�uc�VKa6�?_w�����0Ŋ�o�j��`�W��J]�P���~��"����c���2���<��!}�}U3ڰ+�LpZ��^�����$N�+G�_#Oq	�&
��f�ZL$J�Z���[���S^��[���	Z�h3L�<x�jh��U/%����F�SP����-G�%����<9��~ �쑑>̉e��s�gn�G`W��'-��Kb{R��CrOB��V��q�#�y!k��T��i�`ź7�/ ��6�{yBk����Ӈ���TV�u1r���2�h<�m@@d֤��Ce���erC����Z������;ƣ�Wl�`
L�V?}���ML�y$�P$ 2ԔM�{�+'7
�{:�ܴ���^q�u�Q�s��q��p��4�S��6(~#�
��Q&����O��$�"�J4zS��B�I��	�w7iqNw�S��;���"�Y���)C�x}+�G$%�����WV��������ӿ@��?_H6�}�_���@2�g�5���wR�=�|��/�DB4 �A{~S��ʥ���b9C�K �$:�q�cw߬�&�H�_9ju�Q� s{��^Wyث�%q�:�UL�_�B@"��=ZP�-�F\�u��b~�*3��z��_��ƽ�*�#�������^���X��tc���B�l]M��ɫ.�u1�)��j�4�>�ҥ��JТ�*Cp�}W��G���~5ꍖ���=7٬sŁ��./X�س$0����F��xp�X��\��W��v�<Ҫo�4WT�ܢe�8���ۘw���Wq�c�����0g	��aڙ�-a*�"�%\�M:g:{���n��㑡�vM�w�J㞿�����*���3�)`X��G�b��t���c>�!Mc)�a�>��2�8���$F�iz4����T<yMV�������L�0�m��|�wJ�f87�c�PU��H������mJ�L�	�z��Б�<�ݟm�Z�E����1��.�$�qQ���/��T'O��w�t�]1R�剄v����W�N�H������f��C(rU�a�kྉQ�6�$[�c�tG�R��5���?˯�������N:USB1�VZ���$L'{���H-����0D�O��15�Q��k#��G�@�N'b�skێ<R4��l�a���k��޴�Ո���x�?�$hS��Ţ���L�zm�3q���!f���+���3������eu���dZ J�CH���ظ���z$I��)�Ao
�5F�s��Ȼ|b���5���o����r���(����N�.--���<�f�9�Ȁ��;ķX���c�� h��D���ÌɏWk�3p֘��A���k��s��0_���3�@�WFu��k�y날�-�n�3���d!a)�?�\�x򜱒�q�}��#�<a���<�*�Ֆ�^���7 ��/��yxV��l�7��c#���ᑏ��GL�ڜHD�w��_��'�r�Nld���9�ʗ5���H�̋\������r���\Y�g�1*gj������4�Nm	K<�rR�gbJt�]!�GBj��N�i[(Z�\\�`iLw(�HĨWJSh��C�� |����D�����O�)��+�B��'Y��<Ǐ� ��^�i��;V�'��B� ���^��1v��w�]���;2���W%��T���Of�����j�X4+4B���eBۂ��L��89*���8�ҳ�!��+'E"R1	`Z$穀���v[��X��Ɠ"[�>��|�|)ms3��p�L�D]/{�v W2�S�I����H0����I��''�c�(R��GKp#EN���Jg��a����±'����|����������lXҬY��f��ξ�e}x�Q���*���(�3c�����<yB۸��y_���1�?���HC=�57�E�B��e@����K�����/�2�Y������%�l;;a��[q�!��B�Jm�,J��'ݒ6�`r6Pu�]��#O�^�&�ܸ�h�0ٓXn�Z�f4{�S�p./�Rh���J��8��xHjas�=JM�~�^��iȶp�JL��TI�N5Q�9D�W��K�ck`~O��RK�� O�_��A��Vz"��3���^]%��Z �{P��
@7}�*XX�r�һ�����s���s��ϡ�M$x7���3\Q����y����U?�}�[/���)a��tUW���a�BjL�0D��Ÿe1��7g�ה��:7T�v9m���]l:Q#:���,�c�ő�|��ū�a�bw�;d�ɘ8�c\��yjl���uE�����s�MrJv�u/u0 gqp}l@��5�7|��yQ�]!�a��p��lЛ�n�9~�|DV7�?B��Yn���]峴&����X�<c��m�켰���2���)��k�'�o�)����F�8��Tl�LE�9�9���D��#GeM�A��ҟD���Rjh�-�V�����nr��3�چ��?���K4��� �)i�0Cq�`���r�o�������;(�o� �g�i�4h���*Ԡ�1�^=�U�A=r6����Q:-���}��U�@vi�1VM����8�~��3�,��[�$֭Vҡ�!#��h��s25�L|������!�xIc�D�?�j 0�@#�f#��>��,��-	B3%>�	i�I���5��K�B?d�+����l��0��1+G�j��|�p��� |Ku�����o���a��4v>�x�b ��Us�����+0���0��4�I9\�T&>,���J�(#U怖a��R���
S|�<S�xʝ5������ǡ:��®�b��.��3���<��)R���?5�T�U?콶 ��螉������D�-h�t:�EVu�mu�����,��A���٬5ڷt�2��pc0��&�٘�6/޶����vO��m;_%�i���]˜�5��A��xAݭ�L��LL�n�1���L��L�  �s]�1J�l���z�he���E�8����xD[1�N�a��3�0�ߦB!�Ӽ���ϑ��v��ݽ�p�_5�P;�q*�O�3n0Đ��-��qz'�G�����J=�9o���][�?ݘ�<KEܧ �\4�p�kxJ���:��_�$hj������ F'���&��o�S|Č�wZq���+�pq`�W�� `��i�@N�zQ���K1��b�C%X��tpű��"����E7!Q�Z��3*��dC�rB�O����3�A"��#h+,|�U���2A�H�.���M�=*	���@;���r�3�ʷ���	�ma��y���8B8�݌��Ϫ�y�,�,(k��-���QL/�L�ֿUu'�a4�S��#Y�AQ��M�,�E�����(q��b����Ƈ�W��@xq��?�x��}S1�ď#������P/^#}�.Z�`·#���@�p;h�kU
~X�oG[ᝲ�e��G?��)�$�\�F=���\�{�4�E�;Ai��'Ǥ�5�^ă����C�滴]�LIV�08��hs��[��8��w��4!*㺗�wO�%L�������JFW��Q셹�����m/W#�iNj�����0������e&4��Dl�h�	*&
ǜ�zV����$���Y�n
p��P�����BJ:}����� m�̉QQ�E�QK'��ʱ��Ǧ�|o[��yB����`��'��dK�4߹@�w �^����t�I1��3����9���9oY��-�-�%�K�٦2��CS'����	t���0�6Hc��w�·z�w�֠��+Sh�����e�-�>JT���%�s�0��۪̗뵐����)X�Eo���毐_' OZ�G�ͳ-���?/�KE���^u�˄��I�(�D{UO
`��h{;s}��(���𽜘�&Nq��)W���ͫO���Z�uc��k��1��3j�"�I�����gc���Ǜ,��t�4�E�얌ao�Ú������|z]�a�.�o��H(�Mh���J|[��qcm"��.Q,�e_���o}�
��5*�
w3�h��M�s&Jfĭx~��x��[��[�X ��o�!g��3�V���<̔�  z�w��n�_Mz�.�Ƅ�����g?\C �Yw�@�noL�{JBx4�X��M`�����F�k��3�ov�H�M�?�U�4Ǌ+������*IT�p�i0d6�%F�@�N�r�㵬�]
�E\�mIe�S0]Ɠ��V���8�H��z��`����K~�m��KX+�3�5l6�ǖNdq!����׸���)Sw.�ٳu�J��(����:��|�m�2�����Z�j�;�<�, i�cԜ��ucG��e�9<�&�<� �Ѡ� � /�a� //���� DL�|��&��7�@�>���	��۠$!���1ϧ�BM�5a([R��C}+���Ɯ��O�@��p���h�ݰ���l�
��UEJk�s z7����}֗��ߩ�_7+\┝��S�b�ZxDW�e��3N2�ɢ���Xhy�W�C���s�)��9
|�DϠ䣸��'���e���|��#G�p �\�w�� I�d����t������ �� dÌ6%��]��ص�E/������x����p���44����듛����OV��@V����(�P�d�sJ]I���K�N)�f�H(ُ��
�}~L��:�c��ݻ(}A�ڑk�	{�B;%'�_px`�b�N/_Zy/�9g�p,|hAL�3�8�0�{�4ߞղ�%����|�XgP+��a�ƫ[q.˷iG[ z���e\�E���[��ӸR����3���b������@Z���1�"Qn���0�Q"*-�1�x/�,��@�&�y��*Kll�b�q?FF�K�~l-LdĎ�>`�,f�a#t�7���~����_a}|D,�������W�6#��@���ĭm�Ru6���7���{����z� ��w����ѯ��T̹�"��l�m��!�u"�� X�Ak�����{ 23�Q��f��z�Y��TAg�쫾a��z^Po�C~A�� ǖ��i�4-�	�l6Y��/'u���{��u�2�U�(I1'Z���A��q=��Cy������Ƒ�{�b�y�Ճ���_EiO^�6�&��L��sf
�=N�~�?Y�%
�'��z��E��ϮH�B���ih5c���-"�D��Z���l�80��1�x����wY*p��Smc��e�2vNb'1��n�7�ܫ�8�Q��C�K�}kB�>�ɯ�<jg'� dߨ����j]��]���4�۪
|&��<�b~y4��Vևu�a�G-jT�f�W9���0�H�0q"y�@&��w#��6���$�M*�������[ؠ�x�&�Ё�$��F�j4��[(��)�j�8�H����':;�yY t���=Ԙ}ã	�V$S��"�/��*�k�a�%#.o�s����#V�w��\_�W��ߴ=U���������΢`�(�D�)QsS'x}�
}��~�:ԝ�& k�j���$��+���3I�M\8�>9���K�������3�g�:){�Y$?0�DĔ>�}���Ɔ�bӂ(D��^ȵ��B�
z�II������^��BQ����'$��Zwv4��M�,��N�u�F2ulg'��J�� ��|��L)��<��7#<9�{4c���g~cg�AiDp�Ni^fF�0��� �����tQB'��.W��R�I|�z�&_��5����-z�!�ł�zt�d���FS:D��W�3T�'I���Ү>ʀ;�3P�/\�5��:}�n���g �R-g�����?��Yb@�.�pBp�K��A��I��Y��*D��{����i5�L�>���_��l�%���q���/b��ɉ����[X�Z̯O�D�����r�}B����&�	2�x,�9����� z�H��?�N�M��k%��u2\D�M�֐}�IWǥmkPiL���1Y�B��0knNe؟���LI�8N��~qs̋�)֦t|���>x{��v�k.�2�xGA��۰�ܿ]�_�.�`�E��i~�$�P9�!	QB0]ۊ0�?Gv#����u@D^�6�d�A�~�YpJ��~�Bu� n�lbԼ��wj�'?���`'n�t��?�<�`n�4�eFi,�a³����]2����*#&�{">�9��4�gf|�J��\ʲ��q�{&�5�ɉÝ�"�Ɇ��hK�J���3eh����-
�n+.�K ��S�K�`F����J{T.��d���tȩ�Y(� 4����[4w-m+�cMB^�X{<�	��̼������"mNE�Ӟ�c.g��4͔����;�{cZ��a(O�Nԟ^\o�hi�,�����vPt�X*�{�	V�r"�/��E��8[r�tE 2-_Z5r/� ����3	��Z���h���BE�Ӯ����C����yU
ע}���
X��$��'��v�*��^ͬ~�y�tf�e�"�5�N�$Z�x��_��X�:� �W��pl�DZ_ņ���l��^B�JQ��4Y�t[�c�|�g^�&�/r`��Q@�������OY'�����p���}�\�$�S3�
�����kK���x�zXZe���;��n1��m��p�(`_܎O��;�T�ZX�c�Ҵ	]i^A������F7J۾7-�~-��� f�����S���H���>�����2�=7�[4D"�F��!��m��TY���}!Oږi���o=̼�_[E.��XO����'e�Y�)C���=����8/�l�Y��[g�Q�1��yo�#�)�����$d����A��S0�\���/���܎��E+�(��D��Llb� f"��z�9�?;�tnf��]��ο\�?ŭ�d�ޒr���T��Py�6��G����i�~8������0�fL���j��!{����IC���O�O0I(�����B�ʃ<ʦA��3.�#6��(<BxB���"������q0�8���g,���3�=�� �����BpYV����ش+},:�v��>6�W�wN���ט���`���5XL����,w�����<�}�c(�dNV~ԉ�e��H����x��C �i����I[�E�V�]�۳ 
B"��������'���ѹ�*�2K���,��Ug�'�FB�o����$٩@u�4H�4S /f}ʺ2�V+��4{�6�q2�᳟>�Q�3!Uc 7���f� ���_���]�	7���[��z�f��k�ٗ�Ԛ%$&r��-�;i-���j0T�*�t��v�����d�*�c��H����aQ1��P~�6��)Ͻb4���6����f���������$x9'�Ï5Y[��<�{kf�~w'=xߘn����wDF���� ���g��_T8Kkob�a]7����(�y6��=Ԁ�8��� ��}��{M�Cz�@�wN�A
���t�V	��!��N�<��(K��l�Kvw��#6c����V4��;�a��H�C&,�؅n
��~�]�~�<��(�2ń�}?����4��1��N}�ť1��t��=� |+�8H0J�1�]����֠ᓑ�Fj�}��0M�H@��J�
V�Ӊ`��� c�tj@|�0ɓL��k8�S`��l�$M�]ӳ��?D�z�s�D�v����H��q��(jWP�����Jw#�r���m^N�I���
��Z��Vf�IJ/^>�eHe�ɃC1M�.���N�JKc4� ���3�����.)pnN*�j_����k��;����&m�0v����q	\�W��iQ�}DkX֖,aW��8�P����8yŌ�`����iP%W3�޾#>iy�t�:���~�?�O��5jO4�i�lM��q(���p@l<b���_��!�dd��K*X�F0b�ɕ�އ��+$������?^F�s ��@|��x���6�S=1�7��	���N����s�y�_���D�̴5~4�J҈�H+R��{kq케�Hܡ۷�����N�M�rԿ�ü,#ǉ���]�-�b[�+%��<�ha��cT�B���
��oHdG�p��{�QX)u�����͐�����:��N��<�����n���J]G����d`
�X���%�qg64_v
13o�L9�~�VH�`?�(���&w�(�����o�ػ��h��������e�è,0�]��<г��)k������ٯ,��t���'2�ߔcj�y#�-D������H�_E�r������t��*&hV��4gd_�WS�%��W!���=lY@e���u��SM��Q�:2��
%��Yn�\�yvO�m1��C$��z���b��h�~\ �����=���ad�EX15�,����t�	V8��HƢ�#.���X�H:J����U������	���l������u�Ӧ4���\w㍭�|V��+�Q�s���!FQ��3�276�v8sΞ�W������_�,����[*�Xl'���؋��X7�ذ���u*F�}�.F�fxp��>��Bp��BHhE�z}�-��`�^U����?���)��0�z��J�{q|����Ֆ�ؙ�B���l?_�#�����t���0@���Mx~B���GAN��ϟx�y�dt����D�H:.�{~�J���y�]Z�{�<�^e�HD�_d��|J��.���'�ȃ��Č��ס�����(���W�RRт�~GT^�ǋ�d��>�_���rk��z��/[}6t�*��L��8��I��X�G6�-��Ab �