!������A ;� U�aW�����e�{}�q�m8�~�M�a�rB�M혋d�u���@2.g��_��f�~��:�Ї$���`pF	|݂�� 	
�  �̙�z�Ö��M� �֓>[��\�a#_�R��SY���~�|uԀe���q�Щ��N*��W'j�4��㗟�Cu�By �`B��K=q��v{h��Ҵ�G+�[�����J�9f�U#(� �&0@]P�0���bp\	yW|�,b\��(DL5Pl��4�\mԡ{G,�媤`X�K?�e&6���j����:@��߇IԿ�9���L��9�B���� 4�� �#��/ﴋ&d��un���F�%�$�L+�C$���PT*�(���g��U�������߭���bpy	p�v{<fH�b�l�H���z�R�J�x:ju!�[�@�w�S����#�]-<��A�.8��D3d!��6!������E�t�Fi$`���P��'i�vl����e�O�e[2���жWe=�z�}��� �E%ժk�7 �q@k�x������bp�
ؿv˦  
Y�F{��j��2��3��F�+P�aC���.1%hCs�PM3���fsR�#��Dhp�TW���ܡQ�0�)d� �V�n�uV�qYLu��֪y|��������z��O] ���r(5~�CI$�J�� )������ʵ��`p��z�Ǡ ��u� KH��qU��&������"�O� �A1r�@��z2�D/ͨ	��U�p���� ���X�P-8퍦����t�|V�C<yQ�e��<���r^�Qd�wl֫�C6_[t�t��B7�����6�rX����#�꺰��b`LX/�/� xg_�  w�G�8"ݫ�t��W|��%�ԭ�5�|�=n��?U��ܨYg_��[�bAqu�'4��BG؊�kk�Fz�L"Fw���TH�@%T�
K0��E�d�wK<����tmqޓE�ߑ$0더�J)Pu����|IOcE�t����bpc	 �~�c8pf��FI�����؟�YX�M�%�Q���yÈ�whj�5
s��ݻW\���UR���j#Jh�#�y�P>6A���3��O|�YU�RW�SwE %��U-XU��d��=4�Ο�跄��0�I�� Y�j���q�ے ��`p�
L�zߤ p��YB ���C"�Ɵ�����Cͽ.6j���x��|2SI�犍�)�Y�i��O�L"
$�z�f�n3j*S��;������wI�i����uS����ͥ<�Ӓ�E��H�I��@XSQ�Qy1��1�y�����bp�e|�Ġ ��>�� (2��FXЕW2Z�ԊM��)e*%�3к�j�%�i�tu���.U��q��q8]UR]���6���q[�2#N.I��O��lϨĕ�l�	��[V��|�Q ������贋ɶ�T�`�@�a�襍Py�A�g��bp`	d�~�� �3�  �U?R�=Jvds]e4 Е��`6�c�4�]�Z��a�nBJ���Сc3_�geKɎv
a�Zy�����������}�/��Κo'N�49`���Rv���*f&J �Q������9���4�B�96��U�����bpz
ܽv{<fH�2�pH�q�:���x��NP���R����Ǹ�M��f'ʑG����@j�6�Yw%˱($�<==�bzQ�<��Dqf)!5'��3��-���\D&�����o��J����I����y�@�Ef�� �E�0����h�>k���`p�0�v�<�H@2�p0���G~��7o��=4���b"�$�!`����ӡ!#�	&;�TG�����������wj��]�W(�C�W��]�Q}��6N����f�:=^�:���Y��r���f���,�~��-DK�4[IDuX�
,���bp�
�Yt�<�\Y�l@�qd��������L�fذ�b�:\�O<����vS�g������j������J��Y�d��Q�Bg|��İ6ھ p��d~�k�L�hm��Ǐ⵺�	:$��'/�K���k�k	����=j=nF����bp��v�=\�(b� (FHL���� ��z**��v���er^�'���g�֭o��zwV�(��>�@�#���ڮ������̀E:�'ėe�>���iP+.@�sO ����`f�����\skbD�Y�+��s�[����vH����H���bp�
�etz1\	�z�p0FH��P�>�J�d"��H���_����G@�[)�� �`AbQ��aB����;���.���$[ɩm���첧*�#�����S�1��Y����lI� ��GH����'u5���x����Z�xh� ����ٿެ��``�	4�x{,(HH*��Z�a�Ů&�gd�73�+8J�6����d�}Tn0!��mCQ|D�d�1��ȭI�^�W�h>#������Ww�������e�����±�$Hnu�u\xn�'�vn8G�X��t"��Rq)6�5�g"/����(���Zd��b`�
�tk<fHr��(FJ����~���s��k��O����GS3��~x�S�ˣ����i7���5��X� ڛ���-7��_��ՒL ��3�0q^�@��\��v �j��nU�:��U��[�:ƞ����[s���\gp�	��bp��z�<hZ�1�\Fp�����JW(��*�T�"�jT1/���4�)�t�V�V��ڴ�k��ch1TH�j(�QuZ�a�gLڄ^��D_���?ˊ�h�c"�4m�jW�6�������#9w��t����Lئ���}G���٧����bp�}s~�<e\
�_�H�5��M(l@<q���!A!�e��Q�ȳ%_W])�5��̭����j#�֖VK��R�4J�"�G�/��℔4���P8�R�ü��*��#�T�� �Y��;k,�ʷ5�x�����h�+7�'����^�N���`p�Msxj �\� � @ ��KBo��I�&`�@ȴ�K�]�$ŽY�w{�ӥY�O���������ez7G.䳧J�� i%� 2�b�a �t����R0�Wܡ: �V���QzCU��feH\��%���y}�X�7C��ɞX��4��bp�%uvz<�\H
�l  $R����K �2\��Aä]��"��s�-6�b��m�g�m����s��wt�YX�i4�P����Oox�^��7�n�~���[��T4�Z���g�b�C9�T����;�g�ؔƻm��e��ך����D��'D�����bp��uv�0�\�Z�lH�)��R�"�ТԱ(�M�dt�'�/��Ts�;��Y�|�`u��8��I%YHc�Q�'u�)Y�H4�B�@��&��q"��Q�����``\$���:D:Y�m�
���V���ƣ�(���9���G��	4J��d���r6I��`p�=v�<�\(N� 0�(���O"���.*#����T����~���R�z��ߏ������cZ՞:���XJh�?�֚��L��  	@��4l1����P�������9��ݎe��e�?��b���_����E�X�6��w-*�u������2a�D��bp��p{1(\`N�pIF)u:ǃ�TS"���.7!�l��������K=w�����|a ��+��F	@C�����ʖ�?���a�?�w�Q������@�Z��$���vxr���$%��U#�0'�<Wڳ�K�"�1!IRRBdbPp���bp��Yr�=%\��0�px�����Dی�
U���ip6�+�"�����_Өꉻ蕙ēF .�c.�Y0��ӕ�u����_�~[�CH(����p��F�2m�{�4�n�u�o��s؛cR�]ɭ�%���R��(&�����B��~&���bp���t�0iH	1�l@�qH�4`���2�j;��y�5R����T���W�uO����N�w�'�9`�<�K<�FNa%�qv���,Y1|�X☳a�A@- �Z���	�dÍ$@�W�T>�8�o��肠j9�7x��ԌuHt�m���.a��`p���nk=�\�2�X1�!U�s�EK%��DV��Y�����;�,�1�6�Nׯ�^��*$qK��f� S����9)���Rg�ƍ�;˳���~x��"�U��q�,qcuMKx�ֲb���_�ח�b٫�M��"�7@�BH1Q���bp��gx� �\��"�XH�8�"(��Ø�ζ��i~��IYiϮ���:����N�ID���&�㭸� \3V_���j�����N�E}?%6�