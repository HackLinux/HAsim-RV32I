�������xou��zqbQF9A�����v~������b@Mcv������rbU\�����tnily�����_R\m}����{jVJGa�û������ɮ-2CR_p{{~oMI���ĳ������#  	>���������ؓl\SH9*$3^j��������Ŀ�mGECKS^dgiv��ƴ������}a>4D[nz���������UZgt~zpdUJW������|wz~����{lNWhz�������vbST|����|pknx����~UVcs�������rdTNQr�����������},<ITcy|{nVN���˹������w> E~���������ÏkZNA9@Sd`m���������uchvtylgiq�����y_[Yisv�~|���������aTTWZahknpz���������|uhgYV]ly�����wz}�����yqq�������tlheefhkfr���������{qdTI@<Ng��������òd;IKUZbccabw�������mcnfA1*9Mx����Լ���}yoeXOLFVx|����������uoorkluuoz}����wy�s|�������������pelkkjqp����������}umtlngq}{���������~vwv{x��������xrf_ebhp{����������ue`VSNJMSo������º��sfV;:=COYz����������xdQGOdy}����������sfd]k~���������unprnru���������}{zx~��ssz{{����������zs���~��|�x��r�i�v|�����|��y��|z}{{w�}��������{~ruvmkn�x��������{wsnipb`^ny����������nuoTY][o������������vr~ruw�}ntqy|~����������wuzxusx|{zz{{����������}||{zyx~v�|���{|����x��������||t��z�{mf������|����y��f{z~q�|h��jz�}wq�������n�l\ah��{����j���ev�hqr{��c{���b��~�^�|��m||u��}}�}��n}}���n��f�w�wx�xy����ow�}n��e|��v������rj�z��r�qq�og��u���V��euv�~o�x�L�qy�q�C��ph�`��Q��~�W��f^��W}o��wY��qZ�zrr��i��o�W�|��9��l�|v�A��a��[��<�iS�X�n����d��lI���_G��ijr��rq��g}u�tUz��+���dl��?��'��Q��@�}^�n�vI��@��}@��4�v}vv�P��}W�nP��_~�A��=~�~F�v��W�Im�]e��Dm�v�2�w_�:`��h~w���@W�8n�4�v}�J���Qw�_�w�vW�}P���@�W��'�~�_��o�g�2��f�P�e�m�e}�f�Q�p��M�i�y��q��g�v��|�e����no��Y��y�ia�y�h��~�}m�|�u�|�ng�w�`��x��x�w�~_�vn�v}�v��o~���R��S����a��Y���Y��~o��w~��`��h���~�~w�f}�|��|��{�{�{��t���|�}����g��x���p��o����~���}}}~�~~�xy��yy������~�~v}}}}��u��}�}��}�}��}||��{���{�����|���}�~�~~�~~~~}}���|�������|�}}�~��~~}}�������|��|��}}��}�}�}�}}�|�|��|�|������~~~~~~~~}}}��������������}}~~~~~~~~~~��������������|||}}}}����}�������������{{��|�}}��}��}����}��}�}}�}}}~~~~~�����������||||�}}}~~��������~~}||�����������~~~����������~~}}|������������}~~~~~~~~~}���������}}}~~~���}����zz������~������~~}}����������������}~~~~~~~��������|||||||���������~~~~~�~~�}}}����{{����������~~w~����|����|��}}}��~wo~���~��}}}�}}}}�}}��~~~��~~�~~�~}}}��}}}~�~~���~~�����{{~~~~~{u��������|V|��NN��~nu���z���������{tW}}��u|�������{�y��sz{{|}w�������zz���x�v}�||�}v}�w�x��yr����q��g�n��|���u�|���gg�x��x��o��n�|u����u|��g�p�i�����y��w}|�tsz��c���e����qy��Iq��ypg��n�u���mu���w���qi��qp��w}����u�|��n�g��i����s�z�za���ov��|eu��v������Os�ks�{��r����pp��~h��q�qb�c��ssr�qq�~�}|��{U��mu}�~��a���zr�q�Z�Q~�W��||e|��W��g�Y���G��px�Xo�nf��uuI��u�?uÕ^^v��X�FЭ>xp̈2�Xo�^)�ˌO�m;�ŋ*t���|f}��o5YѮRR���3����Gh���hxp��ph�xY��h�py��Y��Rh��xR`����FQ�ć=K�ȴFK_��R`x��L��X_���^�u��e��]u�]��E�~�p����y��L��gvJ����,��NVm�}�~9���aaa���aS��R�wAw�ȃ=X���`L��Y��RG�ňoK~��JJ���P4f��gQAw��L)ԧpYRL��_=w�Ý8W�å@P���<F���A=��ŇG_���~Af���Wn��}A��o�_R���Rp���Y``���wwK��~��=g���oXA����XW����fow���Y`�����rTT����yS����v@����IO����n4v���@J���^Ee����]m����g~����qy��yy���p��~g_���gXh���BR���YL���hRpx�����a[���jjIi��Lo���|U{����t�������ff����}vv����lU��{Um|��ghx���jz���z����xX~��ue|����n~���pZ����jz�����Zi����Yh�����px�p��xhx����o_o���woo~���xYq���qZi����Yh���hh���xxww�~w����w���~o_o��~_`���pRh����h����hh���~gw~��~}}v}����}n}���}}v}���~w~�~��~~}v��}�����}~wow�������xxxw��������|um||����������~~wo~����}}�����uv}����~w���yyi����yay���`h���wow����gg~���~~w����wwo~����~���}�}nnv���wXp����qZy����pxx���~gg����ww����px���~w~~~��}}u|������|uvv}}}~����~����~www~�����}vvv}����������}}v}}}�����}}}}}��}}~~~������}vvv����|||�����|||||������||||������������||}}}}���~~~~~~}����||������||����}v~����xx��po����~wn}����}}~~��~�~~���wv}����}}}�����|���||}|||��|����������|||||��}}������}}}}}�����}}}}}}����|�����|||||�����}}}}}}~}}��������}}}vv}����~~~���~~w~~����}}}}}}���~~~~���~~~~~��}}}}}}���������}}}v}}�����}}�����||||������}}�~~~~}������}|||||�������~~~~~~~~~���}}}}����|||����}}}~~���~ww~���~~~�����~www~~~��~����}}}}|���������}}vw~������xx����xw~~����}�������{t|���������~~~~~~~~�~~~~~���~~~��~~��~}}}�������������||||�����}}~~����}}}����vv������}�}}����}}}�}}}}}����}}}�����www���xw~�����|u{���ztt�����}v~���xpx����~www����}vvv����~ww����~w~}�����|||���}}}~���xx���xxx���x���~ww~����}}}���u|�|��������||ut�����ttt����|umu����umut����ttt�����vnvw����xyy����xpx����~wow����xpx����yx�ww�v}����uu���ww~����yiqy����xxpx����~ooo���iq�����qqq�����iq�����zrzz���yqqy�����qbr�����{U\�����yyhx����uuu|���|uuu}����pxx�����xx�xx���gow~���x��~w~www��~www~���xhpi����iix���woww����}}v}��}}}����gXgw����x���Yp�����wgg~���}}vn}���~o��~�~����ue|�����{dt����~�xq������bSZ�����mdkz���ztd����aay���zy��xg}����tks����{me}������ppxx����~���~ohx�����qiy����i������~~wfn}�����d[���[CN{���}Wgw~����qi���x��wXv����vPvfw����hhx����o~o���og^���vn}n}����~ww~�w�whx�����yZi����oQ^v���{l\d����mIEv����hLGh���wQXX�����XK�����iab�����yyYp���}n^v���owwh������h__w����~ggo����r[[z�����`GLx����oGG`����sUOd������qpow�������{tu����p`ay�����bMa������ggf����hhp����jN[����qi����~ggw�����nnv���}^X�����pppp����y�qy���o__}����uVeu���w_p�����c\\����aSh�����m]]u���}wo����yiqy��������}vnnv}�����wxxx����~~}v}}}�������}}}vvvv�����}}}}}}}}}�����}}v}}����������||u||������}}}~~~~~�����|u|||����|����~w~~������}�||{{{������}}wwx�����y���~~vu����{{���~xx����{ck{���qqpw����������}gX`�����scs����qpow�����tlt���||}����xxx�����~vvv}�����||����||}}�������~wxx~�~~���}����{��������|||}}}�~��~��~~~~}����|��{{�����|}����x������x~�}������z���|��~����zz�����~}�|��~}}}~~���������{|{{{�yxw}|���������eJKh�����mn~���sjqxv�����yjjjsz{������y����zqiy����}vnfv�����~����x~w~w~}�����vvvv~����������}}}|u||������}}~~~�~~~�����}||||||������~�~~�~~~��}||��{{��|�����qarz����y~�����tsz������xyz�{�����y~}|�{zs~~������~������{{rq~}|{{z������sN?Ew����|t����{jipw}������zkddm}�����{�����sjbq������tltt||�����������xppp����~�~www�~~���~�����}|uu||�����}~�~����||t{z����|�~����z{{z�����}|{zz~��������whbs{����������}mtsy}�������|noq������}����wvu{������~{|�����������zrihw}���������tVDJo����{�����{jiipw�������|e]fv~���������rqiyq�������~~wvvv}}��}�����~ooow~������~~~~~w}}}��������uvv}}�������~~~~~w~�����}||�||�|��|�������}}}v}����~��~~w~~~~}}���������t{u����~~~x���y�x~������{{zz{���|}}~�����z�zy�������{{zzz���������zz���zzyyx~~}��������|eW_~����������yxxwov}������{tluu��~~~�����xxpw~�����}}�}}}}}}}}�����}}}}v}}}���}}����}}}}�|������|||}}}�����~~~~~~�~~}}�������|||||��}}}�������}}}}�||�����|���}}}}�~���~��~~~~}}}}�}}}�������}}�}�}}}}����}~~~~~~~�����~}}}|||�{������|}��~~���~}|||{���������}~��������wwv|��������tle|�~~��������xxow~������||||}}}}~����~���~wo~}����������||||�||�����}}v~~��~�~~~�����}}}}|||������}}�}}�}}}�}�����}}}}}}���}��}}��}}��||||�����||����}}~~~���~~~~~~}�����||||�����~~~~~��~~~}}����|||����|�}}}�}}}���}}������vv}}��������}}}��||||�������}~~~~��~~~~}����{{���������}~~�~~��}||{���������}}vw~���~~���|||||�����}}}~~~~~~~~��������||||||}������~~~~~~~~�����}}�}}}}}����}}}�����}}���|||||��������~~~~~~~~~~~~~�������}}}}}}}}}���������}}}}|||���������}}}}}}}}���������}}ww��~~~���~��}}}}�|�������|||��}}}}���~~���}}}}��}}�����||}}}}����~����~~~~~~~~~~~~~��������}}}����||||||������������}}}}}}}}}}��������}}}��~w���ww~�~�~��}}}�����||||�����}}���}}}��}}}}}����}}�����}}}}}}}����~~~~��}}}}�����}|���|||}���}v}���~~��~~~~~~~���~ww~���}}}���}}}��}}v}���}}���}}������}}}}}���}v~~�~~��}�}}}������}}}}��w~~~~������y���px��w~~����v���v����vv}�����oo~���vv���v}}��~��~~~w���~ww��~ow���wg~��~~w~��~~~~~��~wo����~~��~���~~w~��www~���w~��~~���ow���ww���~wv���vv����uu���}}v}�~o~��xo~��}v|�|{����|m|���y�y���yq����wf}���{d����ww���js���|l���rax����|��|u����gp���ct���et���cc���qhh���_w��~���hq�����yq��qiy���x���o����f}����{l���mmu���wo��y��i��x��w_}��vfv���fW~�����pppw���}v�|��u�����vf�w��x�i����bb����ix����g^���^<����_Y��RY���Y:x���FF���J8�ƫ]@v��vWg�����p�p��h��`h��~_w���xx�����ij���z[���zq�y��pw���n}v��nv}���_o���pYx���>Y���RL���ggg��~_K���gA_�ăFG�ŮY:`��xG`�şBLx��oQo���fJ����^}��nv^�����w�x����wo��}}��]Vu��uDf���oAh���aZ���h`���_P����<W���W=g���`Yy��`��ww���u�]|��m]W���w>����Zaa��yS���Q�~��X_��opx���p>Y��Rww��o��~p���aS����rHy��px�oo~~����yjr���|dt��s��T��po���}����V����}Qo~��YL����Ra���ap���pBĞQQg���n8n��~Q`���yyy����i��Y�o��������l���u��~wh���b��jz���Mh��~o~��F_���pS���j[z����Rx���fv|�u��}��gh���TNr¡ySZ���n}||�l{��ltl����nW���nPn��}Wm���]Du���v�~�Xw���Lh���XQ����gX~��~wg���oXh��gw���~ov���PQ���oY`��hGh���oQw��nP]��uOu��];u��nEP�ÕE8���uDe���nEv��Qw��Lx���:Q���^(O�śNH���]O���QK���R>Y�ӖF8n��|;I|��m;O���g=��h/i��i3B�ߖ55v��}1@���@,^�̇AA�ԟRCi���Sa���Ma����``���K_���oQ~��wwow���xx���aqy��SS���SCa���RGp��x0`��~FFo��g9w���A^�Æ@n���W8v��v<E�æQ=p��yMi���[N���qYx�Ć@e���lH����wKY���bc{��cTr��_g��t\���zkz����^n��ghp��~Qv���mul��uunv���Zj���\d�ËAN���oWu���UGs���VO}��phh��qZy��ow��fVm���NU����Ud���uIe���e]|��vff���~g~�~F_~��oFo���FK~��w_`����La���hp��ggv���W^���Y`���Tb�����bz���LR���oKX���g_o���`h����xp~�~gg���wFw���YRx���`R��A_����ff��vn}���o���h`���xp����hp��iqy���[s����rbr���ph���Wf����me����^n���~gX�����_~��ww���_X���oo~��~_g����w��~~~��ww~��~oo����o_w���~~�ww~���nf���}WW���vP^���v~��gQg���~_~��~g�w���wwwp����h`�����h`x���y����jj�������b[z����pwon���{��l��{����}no��������ii�����gg������n}vn����wg~���xx��xx��hx���``��`p���yi����ii���xx���gg����nv}���vn�~w��px��x��w~���vf^���mm����no~���xxx���ow~���o_w����wh���xiq����q`x���xpx����~~����~pow��~gw����ww~��w~~~����wo�����vn������}�����n}���}v�}v��|�|�����������{t{���|�||�����w~~���xpx���yx���w~��~�}v�}}��}}��~~w~���~www����~w~����yy����zrz���qq���}}����u||��}~~~~���xp���www����ww���xpy����yy��x~���{{���zzz�����|v}���}vv���}u|��|����|}}����ww~���}}��������{�{{��������|||������}}}�����}v}���}}����|�������{{�������}}}}}����}}�����{{{���������}v}����}}������{{{���������}v~���~w~����~}}}|��������{{����|���}}���~w~���}v}����}}����}}}�}}�}�}}����||�����||����{{{���{{����||�����}�~~w~~������yy��������~~~~~~���~~�~~~~~��~~��}}}���|||����}}}��~��~~~~��~~�������~~���||������|��}~~��������~�}}|��������|��}}~���~~~~~~~~~~~~����~~~~~~�����}�}}���}~~~~�������~}}��|{{�����������~~����~~}�������������}}~~~����}}}�|��������||}������}|||�������������}~~������~~����������}~~�������~~}����������}~~��������~~}����������}~~�������~}����������}~~�������~~}�����������~~������~~}�����������}~~��������~~����������}~��������~}}�����������}~~������~~����������}~~���������~~}����~������~~~�~}}�|��������}��~~~~~~~~~��}������������}}~~��������~~��������}~���������~~}�����������}~~�������~~}����������}~~�������~~}����������~~������~~}�����������}~~��������~~�����z����}�����~~~~~~}}}|�����������}~~~~~~~~~}�������������}}~~�������~~�����~~�����~~��������~~}����������}~~��������~~}����������}~~��������~~}����������}~~�������~~}����������~~�������~~}�����������}~~��������~~}���������}~~��������~~}����������~~�~~~}}�����������}}}}~~~~~}���������������||}}~~���������~~}}|����������������}~~~���~~����������}~~���������~~}���������~~�������~~}}���������|��}~~~�~~}����������}}~���������~~}����������}~��������~~}������������}~~��������~~}�����������~~������~~}�����������}~~������~~���������}~��������~~}}����������}~~~�~~~�}}�����������}}~~�����~�����~~~����}~���������~~}�����������}~~�������~~~������������}~���������~~}}�����������~~~~��~}}|����������}}~~�����~~��������{������������������~~~������~~}�����������}~~��������~~}����������}~~�������~~}����������}~~�������~~}����������}~~��������~~}����������}~~��������~~}����������}~~�������~}����������~~�������~~}}������������|}}�~��~~~}}����||��|�}���~~~~}��������}}}~~~~����������~~~}}���������������}}~~���������~~�����~~�����}~��������~~}}������������}~~~~�~~~~���||����������}}~~��������~~�����~~~~~�����~�������~~}}|�����������}�~~~~~~~~~~�����������}}~���������~}���������}~~��������~~}�����������}~~�������~~}�����������}~~��������~~}����������}~�������~~}����������}~~��������~~}����������}~~��������~~}�����������}~~�������~~}�����������}~~���������~~}����������}~~��������~~}����������}~~��������~~}���������}~~��������~~}���������~~�����~~}����������||�}}���~~}}�����������}}~������~~�����~~����}~��������~~}���������~~������~~}����������}~~������~~}����������}~~�������~~}����������}~~��������~~�~~~~����������}}|||����������}~������~~}���������~~������~~}}����������}}~~~~~~~~~�����������}}~~�������~�����~~~~����}~��������~~}���������~~������~~}}���������������}}~~~~�~�~~}�������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          