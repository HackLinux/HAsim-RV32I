�Y�_�v�b�ߋ�ݘ�)~��f�w�Np䚐��؉�U�K�F��|zbFll3���(�+�q�d��YEq��oDj��_ @�\O9���T��Ń�+������P�s��;��t�N�4
`��l��X �g���lp�=�����zM��`�X�0g��T&B����������x�o�/�g���܍O��(���v~��s��� �l�c�~�@�y.���x���hz�&��7���*��￴�V����Ly!8WH�n��CIb�dm]���B�\���BP'ܳ/�i<=��Z�}�z�̐z�{~w�<P(D�(�L�z�OzH| ��e����D"D`f`�u(�CW�HM�đK���"�L���$�|iAi�=�<(�,�Ҫ��$��������8�+��+�Ȼ��!m1�����@���������gP4*,�׶n�����~�`��>���_A�6���@���k�bz��u�`�Z�H(�0苰[���I��ɬ�|�r'L�Tq�F�[���`.�4��'��5�xk��g�7�n>{	��1%?1q �&�B6[E"~y�\�j��X���um���F�m�b�Ic�k\��ʈ�n]��G\&��-���ͪ�z�u���B�N��߆�^#"��4kֿ�(��Ч��G��4(l�ߢ�/@-ZՏ!+�L���$��aYzx��k�Z�[#q���d@O�U���0��Q`��������xZ�sZ{�pe�p���A�q��T�X�i�0^r�����%@�):H��+�Se���;-*��Ls�Ԋ���"�?G���|��Ĥ�%]�5_܄Kd �R;� ;b� K�P,��������x�0�a�Z��ՒW���Z�����D�Ř���E��w�;��gju��1�>�"��'�_��v�q}nsIK��v5;��v�;� �WX�K�$b��sS�����;#�*�G��_�����bx�΃4����h贬!}���F�uÎ�+�����|����y։�dr��u����ec��>�b�ߕa�L	4b��]�˟h\�wا�8dJ�o�[NL?��G�R#>8���'���ݚ�]�Y��I2
����E8E�L��,���Qf�,A�K�P0I�����Mm��y�i��u]�	��=�"��7�&X�'=K����~b1�/�h�=�(��A
�B��k�t W����p�́VW�FɃv�`��ͫ{a��A�����=�`�6=9@�/�l�!s�BM-��Jq�<��A�k��`v4<+E�9�S�5g�3\�r�B�m�/�ׁ_DΣ*�`�bV��a��0�[��*�]q���:����j���<#�2W8娞�:� !#���p�������x��:��gy� �' icN!A��R~-�����ˠ�J^���W�|�` 	����0_���i&��J��2��J�(��:�uM^0��.��J�5ֳT�Q�>p�
�K�z�}A���ef�,y�#	`�0� �.��ƫ�:/0Fu�\Ew:�j��ZJ�p����	;�#�>�$x��֪����c��a ����Ԛ�wٶh��$ ��~ϓ �Dy��z
�Prׇ�g��#���E�Aj[��.�t�~&�y�S�`q�B
� Da��^�̸�2Y	��lZ ���@[
<�r0_Lh��������8� �;�q�4����[�uԺ�ƒ�tҀ(P�N�̄S9\Q����I"��3���uPՉ��&��x�y��f��h]�g�q�EuQ�>՚?S�-���ܚi"�f�R�V�)j^Y�k���D.m ���
dyMM�d�c3�5��ja��Ժw��ՑwAM6�G��&�w<q�����������>{��*U���t�.ȉU�;'YAp����smm :�_;����
f858�QކƆ�{w��k�U��2��&��k�C_G��&� ��,6��%���}�2�;OT	^w����3ϤT��h+!�ȊZW�\M1�$�::(dN$4G�5�!������O����gOn8�B���{�?U��Ē3@obU�x�xk�z�?���3�Z��]�ۛ�@*���|�z��2W�_�3Ӵ����o�#��ؐ��EJ�yT)1�E�;�xP�QB�	#��w�~���MVm������~�g=�_$��$��V�x�_�mw���<Dًv�%j�+�n��X�i����yی�@8օ��*�.7< ��.�;�Ү������7���=%Q^�{�L0�$�"C��d��b��N�~�5�I���c�@�[څ3���L$?�a�ϣ6Za�3�z�E�tN8��Z^���/��}��H��|\N�!>��	<h���@;�Ƅ]'j��3&����ݾ�4��P;b:{��a��O��e�����r����L�-q0�U��_�r�
s�pD��vV~'�0l�I��jE`H"��;���gjMEp�!dn��B��a8�V�{k�����h�a{��J,���}�:4����kWq^�Վs<g=�A9M��l��@(߰˼c����}!/�k��Vh���[l�o��yЮ �ٳ�0=��|f͔�����[g�5FѾQ�u��Ec\|�*]�/;M�������yu	��o��Ӵ��g�E�8���}����c�xA��v��2)׺����Hէ�{r{Gu�el{�g>�5遺o�H�F,�[����#��.�A�Q�M�6�5ĕ��)R�&�=�#�Un� ��_)(�=���+������Y�#Ԣ4Yw���S��H�]���6�aƻ�RNEV���h�t3vjdY��+���3]�Z�]tt�f1��ы�w��Rmc�[����)�n����F�wF=�$g�"�*��+�r�{��ay9	w˥��Nb��LL�ѫ 2)�\��Cu�0tK>3��zw�M�| b�� "b 4  ^ e�o�j�W���wM�[ڼ��j]k��`m�ZS�������vw9ۨ�0���� �*���(��~�I��(�z,� �"����);�  D -��_��X}�>��{{'�/�L��b���ZG��)��]�"T(�e��GNe��i����Dvf�6��V��(� 3P�-}}����@h  d �h
����}����n��F�Xq�؍���@�"`����N�������y��r����qX	E
782Ak�r�H2�q��E�h��+5˂�-Q���!a�D�P$�q�{��m9dv�л�c�]<$@�ID�;��;�`WX�Bh��.�	P��U7�s�����>�f�.�<_�8�A& p<��	��U��ɖ�ʻX�����SӸl���!0�c��ۆ�h�Lp	H7Q'��ﮏ5��ܻ5 fcU,P3�����a!���f�@�� ��axT�*ěBA��(��|��\|�)L�J�@Љ�E�%a&yZZ�EC�b]��d0���A� �(�`�RX"