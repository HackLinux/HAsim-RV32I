X�a$�m��)�.z�퍒�;�W���fR���	�Uz@�}����-�,Wp-t�Pr������%�R?Q,��,���.��\�*�}@��,�l4�=.i"�[<
"��.�j�G�����?�C8�G� r�ꉓ�o;��"�3��pd[q��A�cyv���Z9Vl�bq:�wM�Yp��	�;�<[�F��-f�}q&����q&���2kC%ղ�Z9�m����XD�a�,nZ���,��'>-����)� ,D��ܒ+���+��G<� �
�}Y¸0s�s�o��W�K�k�R����9�+���vC��%�+mv yJ��xa��i�ȉ���5t��˕[k2���Wk�w�h���K��mg�j�g���3(�����Ap�₩R?S�b#��P�����;�o�R��1�S�v�Wz$�)cc�xz���Q$�pU�h6�!W�����O߈�F�y�,��O|1���sN��:T@�v��~�X�2}���,k��]�'W������s�dv�n�n�n~�"���ҩ�;=��SW�4ǅ�ݰH�L�V
�� ��
�Di��QB��O�+�m�����n��X��o��L��4w��G�kԁ��{k��X澓M�	�۷�B���kK����d�X �F%w|����Ym�ЇT[��G�`# �~�k������Nm��=L7.��rm��b���o����3=�r0����٘@�t�_�vp��I�m�6��Q3=_d��X�N_"wr�M���3���%��D'�q��޵᢯z�k�`1"���u�"�2|���}�1��,��vN8�c��	M���4�"+P�����XLL5�,gV�dV��1������+>c�M�Ϫj�%k"�	�J�3�8%�:΋�*�Jr�|(|P�tK��k`%����4����n?h�)eA:��t�� ��[7���)�VЁ' �)��8�?���u`_V;�O44^��!O�[:�Vi��e��Y�#f��q��w�.ՠR烠�:������;^/�������}U��2 �xQ2�pɜR���Xׄk|�.�`�{mSį����0��u��c��P��)����3��:%G��#&� Ȭ"CHB�ṍ����m.w;�p!35OV�����ѕ����n�wk@8�T�H+�1|����7@HҢ�U�iH�D�տ�ȭ�w�{^cuMd��ȥTl��Z�iU1<R����_��X��Z���TMă�γA���~�����bH�B�ք�?U.�>�t�D�GO�'�+��3l�.>�S�j��2tBb~��%霞��=�=. K����RtM5*�2!m�K��� ���lֺ��K3�t"�!�s���CաI����b�|�y��f�,��]f�&����Bk�|w����@bo:��A��㕲d����S���������2�-�/��]Nx���$�]m]�R��k���w1\rV|�r_�WL��m&�?2�<9;#�K��:>�:F�B[U��R[���;�_y틿�4>��]+P�K�Q*��s�N�x���S�M,�ͱ+�ʞ�S-��l4\61 ��n��f	���J޼y�r���dFsF��M�{�c�j�����g���!}�G0H�"o��p��C��o��ܧPi��d�%1�&�Rn�q�q�q����������߷ҷT��q�j�x�xI�D�d��'���3B�<��K�׺�%-6᧯��Fv�^<@�"ߏY'f�"Xӝ�=�"���9�
�n[v��g5�r�rGW�����=c��4��i[Į���B��U���3�Y���vX�Qw$Z���ڬ^�N��_�a�3��I��ۙ�Ŧ%@,�I7�$|j�A�i���t-ǂ�d�_�NMJNb���q�t�}�:�0� K`�)J4�*=)�JP���h�AW%;���`e�W�Ѣ���:Pr����n'Wg�����>���&��|�l�N1t�ƀh�ɴ��	��{|����O o������vf��n���4���s�v=S.��;�^��<�~�!Νȼ�|v�&_r��8Ϧ�;�Η��,_Y3oG��\���P�������2�|�qeh�O��v����Q�	SV��?�~2}��B��	w�t���� �[-�ecfǪ qi%����43�I5��O�m(�q$�4`��E�4?�CWѨTC
>H�ڎ�8���;}��ܮ^��w���.�Ҡ��ҷw���-���ɟS�����3��>6/H*���8��D�C��������W�B�BE�C��\�^Z��F�~��� /�T�"��X�D���R��|�"���ݤ�{u����kM�"��9�J0�.���e�~���!O�2Ed
�T�A:8�H���1���w%�X����IQ+�H��%��:f�����O�<CWw�ՙ��?��K�e~޺zw�-��X<���4p�}x��@g6��kj���WE�l��-��n/j�X��X]U�R����mɌi�N��X��2i�!q��C��Ze���atrέ?e�(C��_���m���3���	��V=�����L�p��pJJ��@*6gbc�Ra�q;/|��Z %��C,�MN�-�}J1�c�;�����5O�s���:�N��1���%�_�y�Τ�0���Q�h���"�`���D���
��`��n���cd-���T����4����M���$A6��k�9E�䤒��Q�V=�=��������a��l�N����R6��֖W���]h!b�YU�w'��}�8O���噖�&?�V����.�WAd�Zi�OjfCfc��?n/��@Mr�&'�C{�jk�^և����»m�L�{n��m�ڧ�].39�s�kc�R�J�l�L<����Q�g3���k��u_xn���`5����|�{���B��h��՘������	�4g2�.o�U��+˓���*'UF)��b+kz�WNq`ZB��'�d�;t[Й����^J+/HRs�qྩ8#�
��i���G��b��70��u�T^�� Y++[ѐV�����;}ȟZ3�]%$��MY���\#'T��C�����w�`/S"g��1ߗ()�\��l����3-$i�W꽌�����ض�kǯ�j��y�i�]��=����gfz�0�:~MPNd�f��KҘ� ��g��x���"�;: �c�o�c2�4����Wr�#��tX5d�."���;���Q�	_ȉ���Vp4W��,��Ű+�������p����gv�� c�c���dz ���]�*e���'��� �Uu� ���^�f<�~���?8�Gu(݃�Z�P<e��GY��s3{[:��������f@��GT�_={�}%m�ê��`���VX��5�?��'�u9Z�*�
��(��_!�8x��c��0"5Sw���l{e
6|�R�����h0���Y-��A}�~�z��t�p/x5��c8���쑑#�~��#]��p"L��z�2��E��#����`W�w��T�4�A����!U� u3R�iݕ�(Rh/G��!�gn\���'l�]���d�5�Fi�YV[u&�=p �L:Me�|�Ŭ�	P3�;�	�H�~2��XT'~w��n*�f�&A�D�Ҫ�����"o_��Ԅ(����o��y�	�x�����/>���_�գ�h�ן�w��`�
vr��=!'%̷o��7	�������1������d���i:�$I�#A�H�t ��8P��3�����n̐*���p��}��,���C��������en���������Z{�6��8���ɇ�G�;Z�5;�^��B��!I�i�1��1DD������ճ�GI�ӷ2����M��w޶;��|����
��o���L*Dݙ%Eq�����{�_��V��B�l~�%��+_q2�2�ƶy��zB���0O��-��r�e�5uu�޻he�C�����pF5����2A�Rj��i��4�s�ưQq�4�EB��f���[,61k�9#u���� F��qUa��55CÁ�i}�~ɸ�-
�1��� �O��/�O��b`}���}u�c��{>Y;qc�]���]�[�HZL/��!zQ��dT�u�}���tSW��P�;�9g���["��rr���y_�[7�)��!U�M� P��˫�E<�r�^�9�W5,����P����d�la��'g-��5�R���s��3�q}�E��odk��Uφ��~~�B+�m�=~��&�#.�Pd=�{�^}�?�����wV��k�m#ԉ6b+�����?-T)�U�X�l���e�Rr������S��$$����ࢼ<�R��['+X'y��So&C6����i���|�z��n_9��g���Y���Z��^������W��a�
?}'a�D2Ɏ1C5D4��$����0P��[�\�m�"}㐢��~�**��=rӬ�]�wWRu*U��܏��B��ܬ_Of��XN�n���{I��c�<�;�)z�͸�kx�� ���6�@�sƂ�	�%_l�I"�J��� �86��*���j$�3�LÏ��tN|]ȉ�9B���{c��6�4���b��쮣�v~&���7�c����6=���R�h�0�8i\1�,IKYDs��t�3���1Cuz�N�گ@�@�r�͍�j���mF�}���ܤ���L=�_f=��W)Q�aʹ?,�ɨMY�O�@:�W��������V�e%	���� G��X����؅L6��f*elӝ4�%A��?�L�1f��,%&�3���Ee��.��(���o�7��R'1.��%['0���*ԓF�������7��j~�Fa�����1G�QjC.�W׈�����RvǼ���_|��g{��ӱ��X9q�^�q5��㫒�װ�ɵ�k<���x��Q�Tn��9�w��qP8)W$=H��>D�������Ǌ}??*^����oQ��g�X�������dZ����R�i���c7g��$&��;T)�O�޿bk��^G�G�[*�dD��b<h�����Ɖ �F���E���0��T���F�y��ƞV�]=�|y�&vI��$Q���+�|֋��P�k�i|��.�4���{>�,k���,��۔���!�I���Et�ГH.��~�ղ�uIQ����\���� ����y�;}]Ys��}[&:��� #|3G��F�uRg��&©/u�����^� 0��^�+�v�?���Ggn�'��S�N��M�:�At��Z��X-?�J������r~�oX[�]�����<s9|�Yg��<��� T����������j�BN��B�mOğ�o堇��:�(�U����7��9˕��ͣm��oE�#�1�ɞ�vldh�vM�@[k�Q�y��'*g������.�r��Ln c:F0/�iz�V}�؍%O�\*;K��A>:ΞL{����O:������)#�׽���xb *s%QN�2j��{���K�g��wfQo`zw0/�Lvo��}���?w �
�V��Q��c�c���@QԮ.��Ml0a�B��_i��~�����at�ZƝ�����GΔ��a�;�!�Q�Jw&�˱������	/]���4�0с,F�51�s)�y�P����(��׈˚e�×RPS�������}	��D�܂��Y�F���!ToB�3e��P#7' ָ�8!h��(�0Y8����	��$��(]r{�����%=
���	ϼ��u����3 
5��c��H��6��[�&At+��h�u��D�8����$~>V��[�ӝ9�L������W��,�a�p|���20�~2'so&#uf
��إ�X3�xN@nĬm�W��n��w���t�Ħ��gqE0Q��p�}�23fܰ�D��UX	�\T���'���O��"�7�I��s����8���:?�o��M��A;=���isB���@���T7�>�*c�;ZAV�ƽ%ԩS�rdaRXI��(;�tD@;_�IP�ab�XAOZZ���U�׈\~߉��#�T���|�����v�C�c�N3f�5��;A���8|��	k�,������E�t.|����4��Cuò��UL��'�}���E��Έb�mv���N`��-� #�m�� ��m5�j|D L,әF}��i��-s�����5m��:�$�C�lZH����Pt2��%��
���,���K_���Gk�k�Jy�%�6�����qk�X�n*A��5ʉ�F`wHeQ��m�2�P��1�"Z,��#Q��FԱ�րg?0@�}�@@�)��I�o�e&8>r%�
����/����ͻ����x�䊣x`҉�K�_k<��z!�k��ć�$�'~���~����Ч-�@��C��t�U��7�������I���H���ۀ�H])����|��o�S�)��'��� ���1ݛ�Oj?Dl�R��~�.���y���dHNx�'�IY3m��D$gKc%���G��0�,s�'��V�=J�Sn��`�GUk�o ����WjI��ű����"B�),r�!�2��U��Ь6����n��g�� A>k���S�_T*Fx�J"ړ�cl�w���Q�wF�"]�_��6IB�䝌�*!�g�C�jы:� �R�N�(1G��YK��>$��U5�a���/&�\�T�8��?M��CD飉z@�j�������*C�Iݵ��y����PW;Ώd��'3�C��ioM`n{
�V
y!�%�V�\@�4�,"�4L2ꖆ4J� A�e�s�@�	��H@g�`��s� ��1�b��E�j��FY�}�Bn��"��&n]@���_��Ԣ�X��쬂���sO��nz�	g�n�^�\�w��1�I���X  ����0l���i,��q}��` ��$�hlPjQ��%������^Rkd�4$��8�zT�ԥ�EN���(����؍я���V��f;\El��
F���@�o %�"�H�����1��\������K�|�ܗ��"��ٱ�R8�q���Z\#���J�ߌ~^P����Y+��c�e>��dh0َ�L}��[�$D�m;��嫊k��!�=6�]s��/���%J����M:,H{3��I��0=Nz'� �Ħ�7����GLB����mߵ;8sx�f���N��^
V�0A�kԱ]D1�T�uq�d�%��ލ΃�h�|�CГ����VcQ�~�Ry<^�����R��V\eQτ6�:�$"x*4���wE��q��Qj����V�g�������J�����f%��ˌBM�8D���HY�6�2F3����ǈ<�~�2\����rE��]a�'�Q=�;!~�NV�^%���)&Q>�V�	 ��xG[%�V�!+'��)�e]�.L�:ʫ��mQ�)|QI@nY��|�Y�F-�_?!1��v������Y.��ڛ�3
=�QF�{��R ���۳�،����８�#,���O;��kO���R_��L7�㔀Z���~�CmN�Ti���v��J����!0\M0\���ݴ��W���W0�^:P[࣐�Ώxq��d!��v����(�vWx�Z����Я3	���C������
^�٩���b�[xN�6�kdXڼӪ�yx�6�l�%Y ��f�Үfdu��XUY����D{Y����Wy�Ex����\�?��(��S=����h{�̒<J�wy�1�٪�0�}�i&(0�yT/��Q�����Wͣ��I��-
7��E���J�V�4p[%&��֞.L��J���s��S�RXYߍs��;�ch?�#g"=��@�Y��E������g�oRI��]%�\ƥ��or�D�C����w��������ּ?��Vó~�7�#��H��ih�̱>q<���RR��9�m�aC����(�t����dՓ٫��0���ur�䧴3x�*T߱��td�69"���kR��`�?x���t���FF�����~�2$��HӍ�:���[m���#�[���Ђ���	&��xW:T�u�ow�NL��(�ǃH�����T)��q�ʰ������A�j
����: �w��4r�B�U�z�����[1P	kƽ�UQ8�~NLpO*��:4)Ẓ謚=���I�cy�%�z xA��a���r��ơ����w���R�x6��3+�����>���ww�1#��I���yj�Σ2;8�鶨��x5V���kO�r�����+:Y�G	�EOV����Ǹq��m�kf4B�std*}��2�����`Ÿ���ύ��#c�6i������m4}�kC)�X��ᯮN�S�]C��T
�:B|]�g�Qۗ�F�q�1�!+p�jT<4����)���Q��c	�F��N��g�1ˑ$*0H� �M�8����.\�4J�g翽��_J����X@�JŐ�6�������Ӆ�Ӱ;4�S+19Z����'��$��ߩ��w<ޑ0<��Y�8n;ס�\����Z|�F�y�ZL�Q�x��a�y6�@��f�z,��Ip_�O|:�Վ�:N���"Ti��RH=�3�#�i6!-p�Z�l�#��R�fC��K���(�L���ǁS�g 3�;7�sr #��ؖ���n5�՟)خ�GS�՘N���2@t"�yK�>���e��$Sx�������>�&S�c�X#�""��źw3|�;���V/��{���`��Sr�t�MW_�r�M�Sh!�������#�_9��eBd��^'jsX��<N�='�u'�k:�/�$,���d���QOO��%�63�A��o�L��Ʈ�*�� /��5�9頧��C�O+�3L~��MÀ�<��[����[+�W�u��Ba�JP�.����[z@Ov�`�k'W��N�o��?�s;���Ƃ!آ�}��kf�fԑ�`R�W��A��s�N����*���Hi�%��2���;�ʵ��e�t���?�"�<$����΂Y�;:uD��z�v��C����hrWn�p[v=5=R�wW�nx�աM�w�9/%����$�ϹT�������[�R2�!�y8�M
�א?W	�$�/_u~A�����L
2��#���U��$_r��(����	}�����8��|jɑDf���k�1`��y���z@t���-���ע�P}}!
�G���@<9a�P~w�C�kG9��p�'��p�q7E�[��ُ��h��1RMx�DLQ��l�m'�,W>�V�:p!hU�����[��'�~`�.�	��4#[�}��������_K�RC���vA�tX�=�h�9�ޣ3���J�OD��k��Z�A�/�8�7�WjvZL�>j���?'o��S>O��v��Wdo?\逳������=�_{����eݪ�E���l>�Bof�:�vysZ�R,��iےW�!���$�i|�l�%�.�?�|"la�Eu� ܛ�yd٪Ė�x��D~Fw��,�3(�D�1���K��+e$�YD��A2�5���jk�2g�,�@���	i�*0�N%FAV���5im\����dR�=9�X�v��E���9�x�r @c����'�LB��.Ǳ�A�M�C�%���� �@Ҥ붪A�#��J�9�0�w�q�͹��m�U1���w,�8�?��D��T�Y
��-�>����G�P�V�IY����H�Xxr)��+�]$�O6JӞ�I��f�򶘸���0�e	ۦ'3;g9�-�C�]t�b��j){��D/%���@�R�M%�`x��-32[��.^�V>1j�Z�=KP�[kr� �F��?���fx�z־�ƽ��������V���*q�3�זՖ��.��^,�n����z�y�y~Pzpz��^�8��X�`-[����TZ��X����^Ϧ)��/��%�����琗�b����X&6�K����<
O�[8|�|�QO-�;w��>|�W�=Xܝ0�]\��P��X�2,3,�̦$�֑�2AZ��C��U�X�ϟ9�j�?�x�1,�f���G�ȄPi���J��V@�- �����f���Gԏ���f�7)5ga����.A��������[5�W;��o߬@|�����, �\�S����ć�W�W:��O�%�ς&E�^�����ř%���{ⳣ��-J��^�\m��Z�^�$���#�|��rx�t��y76b����������������0�ϐo��=vR�}���N���|((����*~&*�;�A�~�Ih��3���!��#V�T�͂7�3�zOP��m������V�\����9�#�m�MUx�mt�%��\�s1L��!��u�u,�T����=�^�c��VT�8
;�I[,�X�^Xϲ"�Q�"�P�.�837R��&;�+-�+Ӳ��k�z@�Ș���ȶd�����������Gj����հ9I��,�YY�e��O�Vu�&���p�K�kU���NfB���k-�ˮ��NC-�}���>{�Ʌ0��c�~��_�$e�������(��N<ն�JrJ<��.6�mL���/F۽�8d�޷�c����>�����*��}j4lZ7�E/zSW˵+�TK�c��J>(>a��[����,m��Nj�G�zx�EÖ��k5��Yy�/e���f[��6��p
f����
5w\t�΢}��**lX�3A�Z�{U�z�F`��I�H�
�"B_=BUV>g,�П��qa'ؔ��LC�������eU� �dmq�8s)�n�|le	�7�s�P�mڷm��$l���f�~�n�0����orH\�;;�p�1���I��=��L��=�r�>jn|��RbP�	{p5�v(r���fS׼��º�V���X+�骊m�;��xث_�׹ ������Gےϼ��[��r�k���3��"�OJ�n+�hsɠ��e��o�]�� 6mk��ϹC�%��{��6�ȥF��9����G�,a�N%w��k�I�Y��+����#�`��G!?0YB��5}K�����g�Ut��v�!��w)5��匍�
�R���2�w�l�oҤ�����J��a�Շ��sU����d�(�9`%dG�JSy&7��)�T����ߐsn��LT���j�_�s�+���bk�u��0�:�n�k�V�B�W����;��YI�t|���Q�c���Ud�Ԩ�Ey̗�[���eH${�3��fR��|{��8ԩڣ��a�U����Y�.�Il�U�(�m��6x ~��;���QJ&�άsy��J_���w�6'&��!��-��Os�9>����˺7c�����6����T��t-t��#����V��}���y��`��	��V#�u��n�n���o@7�F�777!71797�7�7����'5���YKp�x����2�Xc�(�Fҕ&O�j<��,<�M�'3�2�D�&�1�]���=b_�^�^���_�^�^�>�^:_چ���+����{�?�6m{}-�����6�2��>{��*�,]���C����rUF��U����gl����\\+��_���틚������E2؞�y�u+�2�h����ܨG}�Ɍ�1x��֚y��sق,��5>-�\��l��U��l���Djo��F5��FNw�'c�B���g��o*Va��e�,[ҒZ>6���l>�9w[�|�sÌ�_���~3�� W�7��|�Ν#~ڥ!����FV�E�9{=�l_-s��s�oKc�k5˚��e9ᑵ5�Қ�ә�N����!�yYS�W�0(t�HRi�l����Q֒d9pZm8J�m�}Z�`��c^Ө���Y͑�k��t�z賁l��U�bq�f�e��c��Qv�,X۬�b<�w"l(��#�ꦙ��Hugf�U�;ͷ�����4̍�%���;�\��7�a�}5� ��Ov���s��q�h���CVNK5��^x�1s���nXiag������6ٮ��gt	;�'E��V�#AmW��q5Zx/�l�Thl)^�X��u��u�j��T��?_T�,H:yD�9����Y�����,;��~9�8�x�&-��j��8��$nY��|}��9�S\"J��[����߇����}�w��a��o���0��_�LB�"t�	B�+ZWvnv]S�=u~⣒F�W��B!�"�B��ԢE�է���e����ݽ��q5�5��.�Q��3�~<%���NF��SL�h�ZN�\S�`���kgdV9E�zE4 �mh���"B��5<_(�:�{������=N��e����ӇI^`jE�| 5�ҩ:�t���3G�
�<�~��g�ۨ�[μ��cS̐��j�-���G��K�G�i=�/k�#GXc�%��;�1�G�X�}V����4z��bsɅ8i=i&'*4䌥��;��OkVX���G��!���-�
�7嬁�mf��_��VY��K�E��)A��x�Xs���넬(rd��S�ŋ+)C�(@X
-����֘W�j����.�{[�䑋�[�$���)�q�
�����ȩO<�ɪ�5"�0�^2��N���G8�����)�G(�;�ێf/���ٯ
�:<���/���v�\������;�W�ͺ��m�۶m۶m��8;Τc��Όm'�{����:ø�UUO{��� ��r�B�����8E��׭�� ���6�%mc!=�olCv&_����59��'z�cK����;�x���3���-��{��?<^=�_)��(��š��Dh�fd�Q����wl_n]m���y@ً�c@/���`�a��c� d�Wai D��{�:�\L��^�r��p�،�͈�#f�����i�p��
�2����y��]O��F&h`�!���:��ݵ�b��a��O���$?
�%mѽ��8wk�:z�jM
��p��dR��|�|�L(�#^�K���4��6gG��JH���-��XR�v�W��m ��?��i,h��rc<�d;�]��B�*SO�x�pq���]��!z+���[G����3��N�Y�_��í��Pa;��)~Nn�U�ȣ�~�k�?t@S[�ܢ'��߼����g��D��ꔚ�Ҁ&s�e��w�7�P��k���o$���)'�,�v�P���ByN�m�$�c"T����M�a����f�Gk�ݟ3��]�[9p�*E�sZ�[�;�m�+�[0�ۜ�]���ƷBASx��F7܋� 㾓M��	S���X�-l� ���,����Zh��� 6�3΃�2�&
iΑ�Y~���n��̫1��7؋;a��hG
f�wvrW/�����j�+������{��6=�l�ႆ{iX��u8�p10��ߡ����(hJ����o�̴�ZhkU�d��t�U'�?���(d���!����aI�b� Ն��Sң��Ǉ�����,	#��u�ѿyb�i b�"{�T0p�n]Pc㵈{�⇫�J���W̆D�Y�������o
Dn
DX^��vl��mnD1�u�� �uS0��v��w=����P����?6�G����/Bk-8�;�t���r�+����u��<_�����RU._��ه�����>Gbs^:6����3����9��/�C����+�/X��`{����2Z��*6l�4��K���F��e�ڬqS3u�5/Z�J�nI����S����H) ; �?�-��%��,w�v��5�[SN�;hZ����B �S��!�锴�4��jO1�/�������{�IJ���w���N-����[ZY��aG�wΘ������ΞUoox���6�
�G!,ݾ�/sy���(|I��*���wݶ��t�b�ϣ���^�=�Ce��S��1�mo��M�]x�r�mp87O��*D���O�k���mny� qʊ;Ux+mab|PE��RX� P� ��������.���G�Z ���=] �HD�L�\��;�'�|��WM��"n�W�1+���g{2t���eƼ��h|ٷ9B{?�07y��Sٕ����y��h�N�+����D�U&w�BZ�\w��C�Lf��{�
�ď��kZ���r\�f�:
qM~�lMrű�D��@Zk��^�9���0���J�M�� �!��s����:��2�ȮlҲw��$���oo
?�yE��S��άǪ�^��<h6�'$�y�)�,ƶ3-�4ŵ�:P��~#=~4ɒ��&Q�.��a26{<����V�۽8���r�/���0������!�Ev��C����%Ѣ2��~��ݜ<H�p����Ne�Lq�b��Q�O�k,�*c�����J�D�#��v�S�X�����������m�� ��o�A+�n���� 9�&\�3��I6�-Г�$=Y��DD�`�G�_2z_�h��3|=O����9�gT#X�s0lL�
$Ǭ퉗4Q��R�o�>�&9�XY��WW�zy:��o&��1�C;l��� "�a������A�O�%��+��J-o]�}��X�3O�6d!�0n0��?�q��]~�}��BT���,&.�_W�Y��P1�H�{:�ެpx����B⦚��o�lI�C�ʁ4���ZVp��;���(�g6Í�2�2՛b�ᴨ�c|9~��Ar�o�>V�S��(>a4����-�� n�KMY��Q�"�.��_E�c6(+�^yQKw��L%�?��d�~i��]h���"�*���1h��	�&�*a�/�f��QۂP���Ռ�l� J�񭕂ć[K���R�^M�-�A9a�'k�,��E72J��Q��=�,ՠ[Th�g5��֢�r�v�����JӮ�{9y�� ��Ң�?�[���:>��?9)��U�ٵu��M��Tص�#4�ǵYs�ԗ��nP�3�<.�V�pkj��y*|��OUު�+�O̬�k��`�����}]�P=�v�V�K�+�2Z=��tq��&L ���8�	r52=ٕ)��'�y��;PIB��E�&M곡pIIq���TYY��Y/��1�?6�-����e�'":�ȓ��$�He�XI���žMx��N��@=�sG����Ѹ?����a���o.IɄ�4&����V�k�P�l2�'����/�s4��T��Ҟi?�<�8����0e3�qg`2c������F�ׁ��goE8���A�Db��%�DTu#V��s��5X����K�v�u����t��� s�+��V�@&	��Ɉx�ؚ�}��e;�cIK��n���T��9�A����x�{���J�0���K�?������7�3B"�L箣�2�pS!�?=�^�՞�q�]<�N%���eZE%=�<�%�Y��t��Gsp��@h5��JQY��
dW\T3HE� L��8�gq�Q���%'��~C4S�3>�ș8U��7��C���jKQ���\_5Y|e�p��9$M�~6ۛN*��6��Zs=b.��<�2����Y"y�t5s[�a
�g�zL/��>���y0�>M�T���=�f�%�_39:���l�9��tj���<(��e��|�ҐvEkg$58}�E��f7���(;�ċ�P�>v��T�JX#��-M�N�m_���g��*)�C&�a<���������d_x;V��w��s5�n>�i�{0+�ـ_!��x3��唕��c��mi��f��L�����p�2bK��M�>
uǅ��f��@�:� ���Ɣ��f�x��� �Λߍ�	]����c�Rv��ĝm�RȰ�CNO�ς`^��F�9&F�u�c-�EuGQ4��۟}qc&�]h��}'��F?�V���R.Y�4�������7�T�j���#]0b��{S㔚Dد  $�#R�eA��U�	����z�� �vlGb��)�f�S�+��	W�}�r\�;#n��-�y;�4�U�:����-�Ұ��Vg�:uʋ�Tʱ�ը��v55xt�7p������ޘ�{����j�&��%�i��w��9�N��@�m� �����lUK�\�r4#�b����B;��k�V��V��_j7$,�+�o��������~�T]���
P�Yg@����/3��lٶF-���Q2���K� ���M�����,�Q�PWi�|:� ����,C��t���n�6p�^���s{�ˬF��}�=n�'L34�ᓸNprпP�V�Y,�G?!~�i������$`��M�[0R��j���K�n���%��:\�h�bZ拼^z)��a��ۓ�
U`-�(�l��`/��)/I߲nS�wh��d2�������Ƣ�&g�9�bg�=�=�;ױH�멹n��-:'�F�R�`#!�,WIr�)��Y��J���	�_�r;0x��Z��#A�G.���iL�����U���>KRӤ�)�����X}��w�R T�R��O��ɡ�Q�é�(���[r#./�[�  ��A�lDXX�)��J}�/����Vv�H���:�T��ߣj)BC���)���\��]���^1v��9鍿��s��&U�[�8����d$q嫆�t��f�Y^��C=�fcp��Ű�W�~�"�ӓ��#4	����i��;���i��|�0�����Ѣ�O����yU�[�����$�e�����>���۪�:�j$�6���'��}��ß�\1����;p�̋���
C]@�R��#�9�~�� `�����KwZ�4�+��f��{����Xҽ���\�6U����/�>��РN�*'�$��:�
��B��땻*��w�O�S���
�|�/�{�L�3����Ĩ-��98 /�����C�w/��*��o%�]՚�d��T�
x˖Y6~�޺����0��O-��p������)s���G�}E�YM�<�����:a-�Ǐ��^���D�^���~��y��|x�Qק�����*�0�R2-eS\�Z͜��-�;1����I0��k����Lb��K
2�'�É�-t0K9�0��T��������k(_�y�{��s�sF=��<�����`�{њM"B�}\Z0I��'%(OzR@3�E8����e�]�{�DI]{���-������ie7��|'�z�dr�1p/v�������8�
���~²s+�PW�ݭܲt& ��p�a��Q,�������� q���`(��Έ��.l��"�0Wj�i���X�9O�H� �7J�p"9urڍ׸͉�+�+Z��Q�+�ߕ%&�q^̕_�L�m�ԕ�3�^�n���3f3�	�ĕO6��3�{�KJ+J�[ ����ؓF�!�$��Ư�3{l
D�I�Ǥ@�c�ʭ�h_��ټְ�s�늁rQ�a��>����%��JO��E �J#Q:���3C�s��In�do�`�De�sI�hI�6�P]�k���B�g	f�.K7�S+�JlS+&W�N<����g4|�*��6f�*c����2�G,�J�Oi�r�P<g9H�2+�'<�t��w�����>(�$��K��f���'�o����Wfc!|�T#ك���E��-��لCH&Q<���!3"0�p���Vfkޞ�yC��F&jk�a�x33&��>dX���AyLn�4��j�Zb诈�SXM���a�y�Q :$ۖ��V\�ysr��݃_H�i[�WmN-��J�IM�2&�uRz�s���#��Bn���M�kr�t��ۮ��^��Y��fߓ_�A#Ò&%�=,dn�c��	�Ҏ�@!`c�����-�`jҞ�Bi�ˇr �P���h�~�+�?o� t|�����t��� t�:�ݎ;�A��5&�E�ҽ����\������$�|p>��k�A\ռ"�A�'�+�����'~�w�*�@}Q�9�|��L5Lн�fn��!� �_8�xwpᚅ�w��2��wYw������,�H�TR:"_�K����M�7���,]�����ef�p�ܮe�6���얕:&]��g�J�J3���#]lcG�F��빴U��Q�!� /d�;�D�aJ�_����G~:n��&ߨ��nAvQ��5�`��[{�6�[]0T�l\=�F�<IM���)�a�a�p�ˍ�W1�6��u�M�o��k�o��S�%D�s�P�'�n�����{��.��=~Zn��L�˳[��]��	a@��]�_x�,/�'���co�vA�eX�Rh�tw.��Oy ���p&�@�Y~�N�B������W�~��j�+dJH���]����<��=(}J$�����rs<'��Ly�
���k�o"�pG�@� �H��$�<�b�І����c:1d�+O�b�U�s�}c[*a��(�3�'�WѬ�;e:�N{K
_>��u� F`�lo�[�V���mq�L'D�ƒ;�D���O?��d�����;��f�ʆF�_y�����
Q��ǝ�i;R�Q�C�}K���7�o���o�?t�_��w\�t�.9��<�a��� HI��Qvc�'�q���/
'�Cc�����|�����Q -s
!l��k��1�m�/�b�0�B�L=����m�6WS��O<O�V+v�8��ːW�,JW����$YH�iG��q�Q�w�~\�Î��t�����	ҝ���knv��Kg�����W�����}��Pڋ*�@I���f�4����q�28aIf�bo��\������k���?χ�.#k���u����\�KoQԘ���p�7cm������U��'�� ĩ�22Eo.aY����E�С�b�Y{%�"J��/+3�py���6�54[��l��}C,/�z����	�?���nI���፻+���;�^B��ʾ���߉�{T�L_?/�j!
�5��Hb�7�(gT��Ddq�b��]���l�6>GSj�xYB�o�oW�)���W{2�?�v�zZp��͖DL�rު��ѩe���hA�g��D��.�]�GF�f�\ג����C�ac��FW�W���!��&Ҫ�gw�o��\'��u�$��\��B+�F��t�ֆV�F�&���5��ǧ�����'��'�K�jP��ێ'�b޽��U<�p�U�y����{ߑ������G�Kߡ>��GO�:���i�n��{�Ew��^��J������������~����� c��N�ƕy�5��<���#��ad�L#r�)=s�VfO"�<{w�8n�� ���Y����t���̄FB�Y���s:�#���w�nY�9���?�w��k�qj�Yb�Б[���p����?�����z�C��p��z��*�w��)�����\�}��_֟�o�l�Lw5��o
-D��䑅����<ۖb6D �����eZ	/�+�J]���t� �m�4@�a��'ѳ�7�{<ѿm�3�T@��[^��/�k=�uen-5_��RP/�U0k��F#&�Z�Q�
ݪ�8*X������Aa����Ǐ�����`��!AS�]C�/g5W����B%]Uȹ�̒4z�[�w��-�Yo]A�Y�6���P��>L
B	����К`9L�X:�m�4O/��񛣩��w����UHF�i��{b	��o�UI0<|�&�ػ,+M��G�=b�A+�����RI;�\��bi��Fya%�2Ӊ*S$���L��R�5=z��b�lj�N*����#�9I�[���d��l�.]�(�:BlV�(LL�/ԛ�H�3���Ft���]Zr�v���	�h`�T����~g�H-9'���2-]:!��.-G����5��M�����(������7��[�+�y�؀��y�v�q[qn�z]=�yI`���R[T����Vα�
�/B"�Q�D�Fe�UUf}�Az׼]�GU�t�l�y��D~"�\�ǩ��W"_��+�	
H�ԠhFpV�V.�ot��_���L��%��ӊ�@���(C�����M��?��m��Ψ��ٗB�P�\�����-��\�H�>p'/�N�w��va8����]�~UQ8S�4y�0��+���Qt��p�T����N���h22M�Q��>[���J%I�v�ْ�P�>�XѬb�P)�j��0*���@��?$��7}�������l���-K�ןu���G/�Є���ҢʓےB�c����u>:�nl�q�%kǔ��``�������������B�Q�V�s{c˫{��������W�G+��le��4��$3��lD)�u$-F�Ya��O�P�g�[�E�찂J<�B:�$*�nn��J�qn�K$+:�VW<��o����,���	�'n��e������*��9��i�Y��I���-����X�%^;�2��畚��:�P��*��zDo�6���h��(�F�gb��>*2�젨������C�^�_�ѽ*���yJęqwH�����`:��,k� �kE��+�ُE�'8�h
�Þ]a�o~&�Úd�_�;?�u���p����V=��͡�LTԖT:`U˴�-�cneR������	�':!��sS���X��jS��ǡ?ʰI�m�q��[o��$"��X�-�^%���6s�e(���:�`���l���3�#)�b#@�ot�>�φ'������g�Tg�g�%�S(6��Bs�K�qկ�C���� m�<Hh?�nA�����M�����?h����������x�H��#A�WO���$���U����ɪH����9��z�B�ʍIa�D�F#%�DE��CWqZ�hM� I��E�?�7�;����������_,��R��SE|���1{��$)v�r�_�2Z*��}��Кi*Ds*Z�qe{Xb�Ar��5�ZiWh2k����v�S2�Kh��l
p���܅̬��r4 �
:�l
~u_��؉�Y��HXRf;b�5�ZF���Cg�'��(��$�&u��y�.;og�����뉝���);m��EJc���,�����a��+^V�f����ގ���.59HА#2��汳~��]K��q)�^$�*����\�l�2�ȼ8�����便��Z�Y��;��:�{їذ<9it�Q��o\�q�Mj�-d!�`�������
�(8����B=~4�������=��u�;�ax��u�_�E"��z�tz6���fh���<�B�H�0�:�4����,N#�p<cyv�Wz���x��Zżo:C���@����y��:'��e��1p�F�9�yp��*��^?&��:|@���YݻV��!����p��:��&8�}�^�l'��Z�%��P�Tϕ[lk�#� ty��Ry�xiHw !A;���dׅ����0pW^����&�� ���rU��}�$�'�3x��6֩B�O��D<����Z1j������u��AM�%!�S"�O�q����΂T �\Ż��J�dg4!�Qn�5K�9�T��n�'
���<����������]l�s�2�[]�����'<jg<�&���rA˄�븒��t�T_��,Br	{-% � ��,�'Z�h?����?T��]ۑ7}k�n��2Z:�ܣ�{9�]#%KO�)�?�Tc��M�x#��M���Y�Te�x��Rkb�X��)g8��j�C;��1��\��/��z~ߏ�	 ��T6x����NFg�S�o�<��8�>f3zPj'�u��"�oH�߰%B#�"�GS\��ʫ�&ڪXB`��'�R�����"�{�޻jâ^��� �Ѿܥ���\�6��a &�gV��T����������D\��J;͛�dt9��pcθ�x �k+M�ϛ��=`_M�Z�Sm����`U��ft����Yoy{r��a�俒eq�ߊ�=�|�� +)w $E.�ts�,����������1ҵ!
sD��X�p�Lg<T�40RSe2��Ji�`���|4v�`�!�ڷm�%�%��X����q����� 9�yg>/CO�mm����rpD��b�H����:�� \�ܾ�]�Y�lK`vn����삀*� ����)���n�_�ⰁZ;�O�������H �Sn�
��[	ܹ�s��{7�������@'^��r|��)�{5�������e��[a�Q���F����f�uC��Ö�aR�"b}sc;��O�a���zۧ%��K�{���*��h�7ὑ�a���a�R3)P���t��O