�����2��E���U,D�鹨���Yj�\�����{�"��x���=��4��ܪ�qi��Z<Y뾈ɢ�߉�	-���(vE�8�::idD�ndl���4��� D��'�'�lbb�L����3ܔ��Ũ�ٕ��fv� �3�eF�%���~�0���L.���$�vL C����y��L�[k���V����I=�߲ �����N_�=)���Vx��y񢒦ܼ�CE'�S��<c�P�B�H�P�!qU�n�I��֞����_1��Ê��fJ��T�7m"��x	������-����uz������?Ƅ��36O �M,�V]�)6���*-���M��^(�IU�w���N��&�_ ��6}5q��x�ߘ��؟��6ք����<p_!:�S7�ws�[z���^{�!l�~ !�6�y������<d�Y�bT�Z�2`�]�e<��s%Vn,<v8
���@�8��p7�Qs�~�>�BG��{�=����@�j!Xt��l�j�^��)�Ù.�L����b�D�޳�R*j�'��ߵ���ZT��_�<01�4$���p�)��i$@kU�&�v!����d�"�����;3��C˲�Ni �]'���J�����`e�2�>;����.��݃V�qk��}.K�2;����m�W�м �X�)꡸V�B����1���Z�68�8��.ޫ�#��{�?�Q To+U<�����<��=�[2�xZ%9r������	��,��cQ�}i�En	I�I�j4���e=Q;��I��^I�-k�hPLW�˽�1�HW��Ý���"�gS �3S �R�ں4g�YRʽ�͓�m\/�p^�n�����}/n�LQ)�z�,��C��J���������+�e�+�e��|*�{P&�o
}���H���o�j�o~�-]0v]!-���<�o�D%�{��<�NW�H�߶ �r0E�.aO(���J�b����}��~�8���@	��m���p��x��A$���N���aW��h���j���!�>��XP	J�-��O���οd;|�qSw�%Q���ܞqe�5�!�~B H��?�V�
-�T~�b+t���C._��~y̝I�[��(�N���bd���]�P��U���FR1�ƃ�W䷃)g��)9+U�OaB���vө~�F7�+�n|�WX�'+�Ҕ�\+��j���z.B�q�|� ::���J_��E�yx7$w{���ڹ�y�Ձ����8�7��(@h#�X9�e(G�]k�4P�h�R�)�V�����j\
����(N� |�1g��]:�o>V����;�}~� �)�}{�2Ŭ����PQ�^�F+O�3^��=�I��J��ƈ�@-῁�FC[n�5�
�+@�bk��d��4J�$)u��*��<�,eyI��]�pQ��o�-��wx������}�v��+�cs5)
�^�H��uÛdn��AW�4^��M��s�"��/8�c����F���K��zJ�Yi�t�y��0Ⓙ�P1'�R�1����˔�H��c;��=��
��Z3V�?�a*0�JUr�G�l�:�4W��o��dϾ)���jJ9��|p��m&��س�2�����Q*j$"7��`�U�F2�OV���'�ca�Y�+���zB��*�wpPRлNI_�kQ�-?�A`�xV���R�2�@Y���囥���aָ��CGP��1�IH(��K��{V
z2�x5��P��6D�{��rxE���xE�\#0�߱E��=��� �YK���^�be.b�f.M��v#��u�Ĝ�}���C@�b��]UD�?�7�u���GA\����
�`<�	��Ǆ5�1H�E��>W�o)�
�xݧ����g⬙QcҴ���r��&�c�r���zem�d-ۣ�~� ��9��e�릠�8�+E�8�� 's��
Ü�����X{� ���lfD?$�r�{��\�ʔ��\�G/��-��u��-A]!�����Lx�n����g����+��������Zu�(`��U�N]��_�	1`���y�*�yk>�w�:�`�B�*<bM8`E-�{����x�q<Q��{.=>v�� ���u����4*�d����_ԁ��6�J�[<��"���eZr&�3�D�O��Нھ`����k� �X�ND+LS�JW�bC����W � vs��h/ě��/vw.��h& z��rQx+QO#<��50r|<����+�R�n���F� H(/�t�EoG��_����)'ў}�)E�|�����|�B�P
�#�@nCG(�ґ���mp�E��Z�>�N����W0���x����5]�L�R�^h|b��؎��T����K�ý���"מ��f���V0��ý�!�elq7�Y�^}�Xͨ�4��&�.��?[��c�0ѩ|`Lc ���6f�[�Mm9ʙT��{ak��6�&.1��9}s�ZP��|^UOY����z\+Y��qĨ���G<e�����~NT�)�t�©6�P���G\�O����tt��(b���_�%�]�+�����^���w��G��ڷ���R�X�8�"cP%\Z�x1����p�_�p��v#Ƥ�n�\�;#ap�5� ��ǟ(�8���)΃�
QW`}�v2ՠ���������.|����B8��I�{�T����ݷЈ<���p������$cuP���_�"-�5�: 2Q.v��(ˀ��ﱓ+ʔB�+����\���F�!1�&�����h�h�܇��(<�A���-g��N�yn�.���h�C��������=�b2����P�BG}l>����GT��y��n~h�j���K�>d~������K�K6x.�3�t5*%��G�:Ư��|���1��2�K ��"�����5	�i�niI�Ӟ^�41�2x�u�0���% �Ә�S�y���;aF5N�3d>�b���"M]�M�����'��qM���E"&��Ⰵ���4�3��e=e�_�M���y�q}�����"��S�m��:���`J��@%� ���װ��2��h�|�~=���j�W©��;���L ����!�����/NqXq
��!���H��+��F���+�T;Э�*	�]�O�`hr���ݼ������5�El+��3\+�K�J7�}�\�OKxڅf���oB,��&�������H~�� (n��گ+��AcǍz�'��=����t�����=,�D��jf[������>�S���7%�C�S�.�	F{*d����5��݆PA���gY���Tv#!� ��]z�Gn�����&Cd-%�7M!vð��=�ɏ����&0UÝ�L�o���m�Y:�jQ�����=��$�g�t���&V���Q�[|;�Ym/�͇�t<��V�X:����_.>Dܹ�aH�q|���������!�,g����$���jԯaf���
茝f����*/г�a��a"�����Ob�SI����Gx��WḰ���k�"`�=�h�����2ܺ�	u�q�}�Ձm)�ZҼG�������K+��+WiA2mШ��>�G�:S����ω�_F�2�Ty�K���qʍ��/��ʋ��Ůhk=Ƚ�����˙��\�}A��93��?�:�d��
6޺��)�-v��ܓ6�j�F��j�1X4�_ɍ�Dm\�g�-����%�'Ӊ�� Sl%��ky��-���ы��=�%D�|!VÌ��Ĝf^0�Ψ�o6Qu.�$y�f�j�!���բb�ǩ��! P������=6A��R��W��¸�ƚ���d��~ė�NY{�Q���ѹ���Q}�[R��:�����Q�	��7��g��u�g&��1������(�۷]0��U�qʐ�Y�h�)F=��Xd�B�7����9�P��.h�$)M�q!}\쾇�K!+x�:;�h�C�'�P���׶n&�Ѭrqe��s0l螤AA��+Əc|b5���=��)�9�Ù�+')�l��τ_HYf:x��^�y�lT?��S�)H&�M�,$�J��.����K-�
�bp��Zެj�y����p���y�+�Vc.S��S�Tj�יiv�=��v�ǩBe�Ҧӧ�e赭�;�eF��ʴni�����kc�*�;YI՘�J���p��)
��-^��OpX�t���W
�:cP;�4^ZE84O4�^V��w��#~z�T�l�0����0��y�L �x��}��9�v���D��Ϯ٧���Ů�;�T������E�qh�m�ǎ�sՂ����h|-�5Z��g4�I�χY��y��K�+�0��S��2�#��r��X�����a��i@���*8;��A��:�M؁�c7cZ>Q���V�:C��.��!�u�N��U4}�3u��ME� =��6�+���!!k&b��ٺ�,m��-ItH,�7g�b���n O6��!P۟�O���ZQ�O���0I�ש�d׵�G��!Bv`�c��c�ƓV�{��������\M��;_R2V���5�Ƴ������c�8����Lc̍e��eV,����^W��4R�#���5t`�$�|�&�ȃ�g��4��`nǂ����;g����������yӸ50�K�3�|'�0�W7��)&��0kcх�����^��K��
O�X��G/�|�?}��6N�����w�5?��jַM㭻I���� (;&;Ӡ���[vw���K�E���w�g�t��9�|	���y��sgD��RXDFw��V�ҡF� o>]�};����J
Eh� QYn�����#�<K^�~�u3-U��w6q)u�a��H���9e�����g�;�u�k��n�V��@u�lBP` ������?�\����=���H��4k�M�%F�_�2q�VDh}�J�ɮ��~�)Ո���T��{���3�|�@=Uǖ����o��ͤ"����߭��s+�=v��pY�[�?�J ����G%"��ٝ�u!�Q΢l��+�����rK@s�*�_�8��
O�?�֛���	����Hjl�IXk�a!i�p8w� \�K�6
w+�W�8;��v�t|õN�q�F&ȪB�V�ړ�s�""���gL�o'~ �թ}�Z���L�B �M�;"�&���!<�q�`��#"#p
gӛ������0��8���TRK�/��U����}޾�t+��2�ο��wm򚏩<աL�-�{U�q>���{�S6Ȟ$�ۏq�B�������_�����
�ZL#BM�яK��G�0cR�a�zɉ38�&�|D�B���#�.BZ�����������|.�Z�u'��OD��b�F���;�4�n�E��w�'VK��W�����|!D��yp|l5��5["l���\�Ҫ��|~��MI;d,�-L>��������C��ފ`b���C���Y�g���_9�����4-E4�杒�6~��9F��W�9�j���W+�"42�ɍwa#k!6X��/�>��=O~&����.ጧ�<�����gW,\B߃j��R90� �Zb���{���*m��5^$�Xo���W����y��jw��-�nKZ�6��@��jp��B[��
�3��>eIk�:|�[Sv��E6��>���e�E�
k�U5�Ȗ�L�Dn���t����2�ҙ	O�JΓc3'vH��F�d�\#�MDg+��(y�4땨h���!U�a��0�����&��Sx�o��GN!����{��'c&�`2,^1[��/dXoP%��`�c�D�D���N�p�e��&�'���ϖi�(�]'�n5Ɩ�����
T�4�&T�9�+��
a-��I�-XC�� �4�"�"�Lo^�U��8U��'Xw�Յ�g�`	���d͗W`���������?s��ܔ8��3 �$�%0���,(���.�>H>#�����ò��%��'!B^�Q�6M1�Xʩ��)w��aM����@{|�6fj�+Ѐ��vJ��]��pW�����O4m!�^��J���l>�xe�/����y�BU�^Qk"�rąe7Q��K.s1��x�V{�OnaЊ�H�G��hA�9Ua���X�T<�I�0 �R�A�W�G+Z&֋Ċ�&v����q^�=L��x�ab GL7#�Xe �Kx�ֵ3^9��j��Ȥ�U徸�Δ�I�0��~Ε}�'bH<S�
�9e�c("O8��������W�z���`}��[��3g�/ӷ�Q�wh�u�_�x�ɾ�@�q%���-@����yQ�M�c���3D)A���N��.�9\���v�x��/@f3�{���~["�W��=�yN���f49�/讍k���L�����.�Iv�.��Q����8|���r�B��J�/��&�x��^m��ˈ�Ϡ��Ubg�u�^������6[O��H�S�K��d�w�] q��Kp�gp�ɘ��O���?2c �,I@d=qU���`���.�,�
J�"G�ԡ~l�L��6	�=j�|Z�t]������J�93�]7C<�c���w65�Z�
4ȡ$1�����To",�V �\&���5��;)c�YzS5��J$�򙽺��!f��L!�����7��D!�Q��nFѽz�s��l��11��P��[���w;����X�v
�6�[�l�Иߤ�#;��"�I�?�}zN'�|�����j�VFxi���=��%g� �{������=���c�R�:%<�n�M�F�"{245a��I�Q¦��γ晻FW��\�v��U>�C�q�Q�'��h�,��D,���Ҙ�a��e6�� �B��{��s%י�\C8v�Q��p*��P��p}�XV�p��"���d�I����D��2��:��