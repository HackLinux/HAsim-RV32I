?M34=� ]#)"����O4'���-�|5N帟&�\���~v��K_����v�;\��y�ɾJ��%���J<�-<��-L�d@'�L�ՂH����Q��և���3Y\u����Y�-;>yڳ?h��#MGV=|��q)A��f�&����^�������d2���v�5��i5u�EVN�Dі�����Oc(iE������D��Y���v��E��ý�C�-�r���Z����Q�>�+����C��(6�e4���8� ��j9[�uթ!�Ծic(!��b3��v!��>�ϭN"��=�׳"���Ӫ��h�MQ^��6g�8%���n"gb��sy�Y��\n6�"`G#!R�^���H�(�2�oW�~�� �NcvG�T�$���=��lG�U����߫�@�����jc��uwm�����d�8��)i�<�ſ
�J�j-Q;á�9���q4��~�2�|���k=�[.�V�&�5�V�LƯ���$b�tf�>�S[Õ7�0�W�?�{x�d�j��Y�M^��k�Ho�ɛ����ŝW?��q�Ź}�ȝ����d�(BR󞠃1���?ƕ�\����������7?Z<�1�)��~��2!&5u��NP���X������R�$�c;6�($��j/���O���h�I��r�ŃWB����Nѻ5�O�Ze1���N��lyc7s<�R?V������_	l�T;hf᳇���ӏ�d�Vb0ш"��N�τ!�s�S�T�H4�w��t�0���Hv�5�c���'ANp	YgEW��:��a�8Z�IL/hJT���m���CSЅ7˷Q*�zؠ���B��EC0�01�q5L����pG����-�ء�(��V��$�;��uJeX��<�_���o	�%T-*����}�����z£:�c���&�*�����} ��b�$&���D'���q!n�-�lr�e������|60�e��S=h#���O��*����e���(��������sڭ.-�K� ���fk��Ӕvw�si�C+b.�G���k��w����-��k�_B���$I��^�uJ)�N���9	A����fJ���?N3��������@�p�_O8�6ȉ��i��|B��i�B�T6<Ր3B�����J�	]>qe�>��!\�%f�vXN#������c	�.}�.+��{���Z���� �3� �*��Vs=.g��ٔ�}��ҙ��0��L������/��Pp�m88��U#'+R6]==�/t���+�RQz�iq��$*��]��J���	t�r��i�.u{E���B��3������2�0�m�75��]AD{<�������������ٸ17��\6���&�DF96�Q���2�,-��H@`���/�L$�rM&��68�ڙ0������a�ݟk�?Z�3����D��[S����9ׁN���H��+�O����"��6	�,'<Hة��V���1����#�����������J}�Y]H��G���A�ܽ���}Uu�)����I��o �$0���ApA�χ�lO-d�I��Bu���i4~�d'R�j����Y?�-r�M�-KHAvI;�b2qcTh�L�Ʊ ���^���I��a�d���~x�J��"sI���|6���J"����y�'����T?@$,��A�qjԈ'Hv����T諗o�/"��
{Q铀��bћti��W��ͭ���!�R����� �\�-S6s�U>M��:.��x'~y�5�"�sV�y��Ȋ�����CCC�WK'��x��X����#�V�H��=	׷hU�x�����w복�,si��׭��M��{Ψ$ݡ�˯�gӂ�� !�da���Z c��As�\��
����ݹ�+�i㇊]�U9uY]��M�MIA��|q8c�m���dQZ=�:�HE: 3���ٍ������D` ^z�7�5�pU����]�B!�ǂ`~�pL�;�W�5�������)�3Yp���H f�562_1?���/h���3Z��;I��yT�،�~F��W��%,�r�"a)�ҠIG��Q�{GFq�)��x��xap9Z�j�i�>���*O�Dp�@$�%`6���(��4"�e�#��%w{ (�W~[.���>��>Z�/�^C3���Oh�P��Q�@�!֕�Cv%��ǵ{Tl؉%|��
HdJ��$���i���Zm�M��nu爚�p����!�#�o죚p&y����I �,_xq���B A�B�H`i9D�C /���X����o�[�ſ�Q�Kx�
x�����z����(vڨEW�/7ɐ�KY�B��E5#�� ��NRi?<��I��N�$0-�y�������`��~$�r���.�Oy�'۴E�^��yχ�a\>���m9�4�j�pYe�W;� 5n��7�*�Ӵ&Y{}�{�'�QRu�um�$��@Y��N�pE�`*���򊺕�o�b��`�<��Ц��07��S)R����g �'�L9!B�M�Lpt9�f��
��}�Mu�fˠ�v��1�JCGÖo:�����`>�#8��&r��[Du���?�g��������K�D�v0�����v�8T��y�z�|�W�g�@Չ����\,ԓ�]��(o�.b)9ٲ-��:��o=���˟�i|�;m:�ǣn��,i��=����d�3��oeq�;!I
��������Kc�BW��ad��W�dz፵܍����;�8�r�B`p��乢��4�Q�^M���n�Wf���B@�Ԥ��³�O�.���	�B\+0�n�����an�}_m�1�E7�4U�%7�y�}3� Zڼ�tm�,���2۫'"3�� a��G|�!=�Hؤ��d�=��2�c1�̭r(��Ͽ�m9�T&������U �e!�5e�K��U_���&�+�ޕIYT|����<�u�r>�L"%�;%K�Xn+;�̝��������sL\/M��#��-I��- �M�'�BUo��OX�SL!�Lc'��pF�X�5;2)=�k�N���"� ��&u�Xgo���jJ��c��m��\�$s�_5���$���#���b0����q�A��)�u�U���ȩ���`;a���S��H�ǽ��45D�b  ��e���d�/�#�b����<<�z����D~�e�:)��O��]���_P�T3/�#��z�b��,�%�s���tH�l����_V�S&
����Ќ]�Tb#��b�N���r����<��Y�"��������V�R�:�䘅������;���^�dv/�#�1���:8���/� �bO�Tk���o _��XP�U"#�T�S����;=��YQ�U��������`��U�����������o^W�S���n�j2�n�R����i�<�$�%�����\�U����c�-���.7���/8��䈪���t���"W)�%�5����q�	႔��O���!���[弳� ��	~�e��������$3仡e��Ra���Et�d�����b�*���l����YP�U"#�T)����