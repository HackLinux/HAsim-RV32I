}YJ�[A�]KidD(gQ�k0lir/(u�v2� $�N�Q=�SD�T&�W?�X3N\Cb>b4�b4�c5?e;pe<�e	g'eg5�v(w68�4M�;P�8Θ<�0�vw�2 'N9-N)O0�O9S3WS6pS?Y�^�e6�e2,g-�l@wm;�s)�v1�1�8��5\O5�Q/�[�[A�^'_Fb8gLbk3FmLGr@�tP{C�|9o�'c�Nh�S����+)�F �ݔU\�Wi�K��7�c�~W[�Qt1 63 G5 @N Q$, N>	N4N?NI$NE-NK;NK�ND�N@OYSOQeQUkQJmQH�QI�QT�QERoR2�RGAS9WS6kS9�S6�SGT>FUM�VM�VY/Y3Y9'YI4YQeYL�[ZE\S�_4;`�bW�cP?e?�eSof@ gJegCDj[fkO�kW�sT�v4�y;zO,{K�~W�~N�)W�E"�D8�E��Nۏ/�7�8F�Vh�^b�?��L��*{�/ؚQ$�L[W4�[%Kb$eh$!\O&OS[W.�`b�5�)YO	sY Rq_ �b�~;N*�N�P]�RP�VY!;`�y��K"�A8�Nߘ=��&`Snc��1 C2 G8 P$
N>NHN-NJ:NF;N?_NJ�N5�NU\OC�OF�OJ�O:ZPH�SM�T#�V=(WG�X.�XG'Y0f[C\?�]E1_Q:_5@bHMbLbQ�cGdG�eL�eN�e5f</f@>f0nfO	g6egM�v�v7zzL�z.I{I��G��Up�@�F��9��Aŏ=ȏTۏ:�L��Eϑ)���Q�FE�:K�G�$">N:�NO0�O*lQsQ=�S4�S'Y(}Y1U\:�_7@b:�e+:g;t$��7w�3l�+�-�R&+Y��&�
NT�NWeQR[)R'Y.�] �]4:_�_S�_#o`E�b9egU�l@2mT�mPyrT�vK�vG�x]s|R'}/�~O��_��a�Uw�Z�5̑Z�dOW|QeOSpS 'Y?�Y�[q�]o;`H;mV�y3J��D�y�2b�~�k'�qN<\O"�R-T8XT$a?Kb;i fk#+oir(u';ua�5��<f�-��-b>�kt�'�R U\�_�e	R�&O@�RJ�R+�RTU�W@�]�_C�b?9e6YeK!jl=T�T�L�R�_/�e7p�4pQg�g!n�$�XYe'h�*�!�z_�l���[�cLuƖ�N(oR1(W+�]�я1�~�RDOS:�V54Y=�_F�b�c.:g:�yGň��Yr$�T@�Y f[�]�v$�wD�~#��{�J�;�N�RC'YCZ9�[M�[C�e�g-�iLmPwm4dq<1r+�u-�~I�J��C�Hf�?��M�O�T�.yQ� 9$'NA;N9�N2�QA�Q0oR5�W'Y7�[;;`�k.�v%�@c�,�5	�:��O �;��;��0ؚ;A�@$E�OY�OL�R0�SVX@'Y1f[^1K`\�b@9eENmWu(uH�u�y&M|WÀS��Ho���\b�&��I N8N@NC	N:*N8]N@�N-�N;MOMYO>sOkQ8mQA�QL�Q&RTBhTB�V9�WIY*'Y	�[HJ\Ht^1�^P:_4@bNg3pg=wON,YO'R.CS'�S/T4�[%t^�e0~v&1 <h*N�X%�[6�[	\8r^4t^$pe�k&$N--N@:N6�N�ND�NC�O�OS�QOS(WS,�T<FU2(W:ZJ\/U_0�cEYeJ�e3vfC�m>
n\�n2yrL�sK�sR5uAI{<�~@T�E��S��1*�Hz�C��/h�AԈ,ڋCދI�3��Q3�C3�M5�O\O0�R$T5�TFU�["T�D���FF�	g���N:7b@Sb)�e
�f&:g4�r�~7��$y�)hQ%�~�NE�N+[OQIQK�R*S!WSG'Y<�[H�[5�[Q\Q�\Q�_N�bP�eD�e�g%�kQ4lB�l;mOwm#�mVyr8�sW�u7�zE*�F܃Qf�8��O�G�!�Cr�V^�2�6N(�X'Y)�[*_1i_1�eC�gDir{v<(�:ȉ�Q1 1$(N0nc&	g~v$,{4���(�e	�hnm_t+�t#��	�OD�QI�V9�X5�b.fogXtmOuo�R�SƉH�A�$*6R/7R<\�^�g,�z3,{�/ދIa���%�/�[:g
�/�-N7O&\ N)(W!�[/�b<1 %2 ,$ N)eQ�p�v"ؚ,$	�W"��*�R*FU�[�w&R�,�t1 W�N �NE�RS�SJ\.t^<�e>g?eg$!k<uDz?�~Ji�E�R)�N6HQ=RR.US+JT=�Y5P["�[B�eA/fF	g.,g;Pg>�ldq4Hr<�tIň$��>'�R{�H��V� ^z�$N5�SC'T@�]Kt^ _D�b4�e:�v5w1�E��*��AۏC�*$�N2�N�S.�W4�WC�Y.^(�~Ǒ9$DN�NOO5�R	U\+b>T�N.���%[�b�; NN9:N?�ND�N<>PJHQ@�Q8)RF6RE�S'T>T1(W,�X;�X:YAY=:YE�[;�[?\1�^@ _2b7cA�cF�c9�eC/f$	gckA>mC�mH�v=xE~{1�J��5ΏBۏ>��9b�>��Gf�1 H N=
NBNIN&N*$N--N,�N+
OF�O:hQ7vQ�RFS3WSApSI�SH�S3T4hT=�V&�XIYCeYO�[=�]G�_CaKbD�bKte?�eC�e8�e5	g4,g?egM'k$�lF�lPwm8/n+�oA1rL^tN�vKw9�yP�;T�<�@w�D��K�7��G�J?�B^�@�H��,�0�N)R[OS7�WR}Y
�#��7�N(�YGSb+�b	�e&����/M�.N,>P!wPGtQ#�R=NS$kSL�S6�W7�[�[?^DP`!b4XbB?e6�k(�l?m>�rK�uE�v>�xV�y6P�"r�Ne�=��=*�2+�?p�6��'��GўI�K1 \2 VD G$5�N_OV�Q+�R$�SX.UI�V]�WN\1U\^2�_[lbL%c1�cT9e?>eEf'egFwm^�s%u5u/�uGhyKh�  �+�^'�Ow�2��B�Xu�[��Up�TB�#�S�N0of@�fB4l=�m�~:-܀=��D�-N:�N@�N@$O,0R�[�[�c-Ye5�e'"k1~p!t-�v(��1Ǐ5:NS�S0'`)b�l4i�(��.�)R�S$sT&4Y+�\
4t3T� ы2�'D�(�fNR�N/�N=�NxQ�RU�SQ�W8TXH�X;�]J�]7^S�^3bC�e4�eG�fL	gQQgQ�gOiP�sP�sF�sX4tF�tGu7;uOxQ]{?M|0�#
�Sc�@ň=��N׋=݋J�Df�H��5��J��DG�Fv�9ΘK�AQ�P N$N"YAQ:iR1`S2�S@TD(W5�[=b?�cGdA/f 	g>m5(u2����$ۏA$qQ)�Tg�~*�$U&�V  _Ɩ)NNK�N�OB�OBPI�Q7)RE�S*�S@TI(W5�[D _A�bIcg/9hG>mJ1r.�yK�@���G�:`�?�G�R%SOSJFUH[Wbq\R�]U/nY~nt'xMT�$ހLD�TΘJ$
N#N<9N9fN-�NDKQ5�Q3RCMR&�V=�V:'Y1f[�[.Ye6�e5�e7�v)x"?z3M|6>(��=׋4\�5��9>m�$:N�S 9e/}l'�y�{)�N@:g)�l zzJ�C��N�N)�vQ)'�$�1 ]NU*N2-NZ;N?�NXOYOZSOa�O[DQTZQNlQV�Q^�QQRY;SZ�Si�SM�SUFUV�W@'Yf[T�[T�[K�[g\NB\W�]A�]]�^e _XbN�bb�bY?eI�eX�e;�e[�e	g@:gEag>!kcl2}l]�lY>mOwmT/n`2ub5uQLu,w!{|2�~%�~[�C*�Mz�f��Z��`	�\�I��c��Y��R �d6�Ny�=��C{�`ؚG�	�\@�mA�;N�ZO@OGOHOB\OlQF�R?T'1U6FU'YQ\Fv^>�^Db8ybQ�bB<h?�l,mWAm:t8�|Y�~N�~W��Q��G܃J%�(D���S�N'R*)R)'Y1\"<\$^)nf*�g	�h.8l5�s8�4�* �
3 [ NA	NF
NGN2NAN1-N.:N?LNR_NY�N6�NW�N=�NN�NQ�ND
O9MOO�O6KQOmQQvQ7)RRMRR�RHS@SHWS:pSD�SL�SF�SP�SX�SBTB	TZTUhT=|TN}TZ�TE�VR�VD(WK�WNTXW^XY�XRYAYBeYTf[3�[L�[T\^^\3�]?^Z^Xt^K^J�^?�_K�_N�_)'`@a!$ad@bS�b;idXteT�eS�eV�eJ�eA�e-/fE	gNgFg2,gW�gZ7h7'k+ek8�lV�lE�lN�lZNmTwmD�oX1rY�rJ}vS�v:�yT,{PI{B{|"�~S�;T�Eހ(~�[ςK�Kw�Ya�W��Y�2��S�S��Sُ5��N̑M?�>^�6�N��Wl�O��7A�$):N7IN;�NS�N+O-R!gROoRH;SBUS9�SR�SS�TE�W8�XJ�Z@W[1�[3\q\;^L^K�^UKbAbX9eJYeI�eM�eOfT�f:�gV!h-ehU!j@LkJ�pJLryr?�rU�tW;u@�v<�vLxT&{P�J܀7�V��N6�7܃?W�9��B͋@�Z5�Ff�KR�0�Al�O4 I$N9-ND:NH>NC_NC�NF�NH�N<�N=OA�OOHQH�Q>RIMRBkS7�SH�SI�S=�S@�SK�SWTJTA�TG(W3Y=YF�[H�[H�[@\/1\:�\DbA�bK�c.�eF�fL gCyrJ�v �zE,{1�~I�~>��F�M�N��AԈN��=�Bw�Jl�)ۏE��C��;$�BQ�F1 BN-N?-N*LN7_NL�N?�N,
O"UOA�O6ZQIhQ=vQ8�QCR9)RM+RI�R:SLSSS>WS4ZSSbSApS:�SD�S@�S?�SB�S-TH	TD�T@�TF�U=�V5W>(WH-WWfW<�W9TXL^X=�XGY<YB_[I�[N�[3�[C<\;�]J�],^@^D�^HaL�bFid?�eF�e5g0,gKeg8�g5<hD'k2�kD�lB�l3�lJ%m@wm1�oN�sF�tM>yA�y6�y?wzN�zH�zK,{H"}<�~=�~LCWL�0T�.��:ς;��;�C(�F��A�3�>�E8�F^�@��>ُAёM��O?�,^�;�Al�4ΞH�A*mlp�$$;N�S4�X.�c9�v ѐ7v^�Q	��$�N,O0R"�R�S!�R(u��$eh
�{�S4_6e�k"�p�~.bSl$��s

N,hQ-+Rɋ�] $
R";m)2u-��ΐ5$?QAS%X0�v�|S��ST�T0$U4�N(TЏ�T 1 J2 W3 `4 _6 d7 b$N ND
NJNXN/N2$N'-N+9NE;N_LN?MNf_NV�Nh�N9�NY�N0�NU�Ng�N9
O9OhOn�Oh�O*�OPP]:PiKQMZQ]hQ>vQ/�Q`�QW�Qf�Qf�Q[�QERgRqRZ)RNMRL�R/SYSNS7:S_WS8bSTpS0sSg�S\�ST�Sa�SQ�Sb�SX�SF�Sh�SO�SCT=	TLTb4TfhTY�TD�TR�UZ�Vf�V0WE#Wg(WXfWZ�WBTXR^XQ�Xg�XCYEYR'YS)Yb*YieYH�YU_[a�[[�[E�[R�[j�[X�[_\Y<\J�]4^`^_^N^qs^^R1_g:_fS_V�_/a4bKbd@b\�bB*cKwcR�ckidOEegteN�eQ�ef�eG�e;�e&zfN gX	gIgcg5,gJeg^�gf�gP8hi<hX'k%�kB�k]lO�lI�lg�l/�lC�lD%mZYmjwmI�mE)ni/nH�o91r@Yrdyr_�rh�rU�s_Ytk^t;�ti1u`}vK�v[wGfwO�wY4xdVy`�yf�yH�yO�ynFz]wzR�zQ�zW,{M�~R�~_�~_�~^MpWI�+�LT�?��U�O��NςB�*w�?��b�Ha�I��I��a�0��W�l�\�Z�g5�d8�\^�\d�Yt�s��=�hُXۏY܏j��\�]̑h?�8^�7�8��d��;l�>{�jΞ\ў[�]�.�cC�9aU�U!� $*s 3��`�u"\5Lr�y (�)ԞG[O	�R6�R;\�g4yr8�v<W?(� ̑)��.�^gR6q�N*&O�T&�^4Sb�c9�e1yr/$*N�N!	g̑�U �N0f[ �]N.�N$�N	�[q\g�N�Q�SThy"�| N 	g9\O/�S+b,�l-8n2Gr$ANYN�N�NPO �QZ�RO�RhT[�T:WD�W:'YKf[A�[<�[:�]@�^?�`I�b/�eO:gPh)�h4�lS(uALu.>y=�yUT�K9�;��A�K8�8>�UϑKb�ZޘU9�R$�k6Vy9R� �e��$fU�e��>kgR�[(�m-Ώ"i_�!Ǐl		T3�[�[�_�v;u��~$�T $�[�3�b�r *N(�N@sOOlQCR$S-AS�TP�V/�WEY;'Y�[2�]t^9:_@bB@bF/eB�e*hK}lP�lK~v;wB�~=�~BT�K��;��G�Hb�&0R�V�['�^66e/�eeg	�N6
O:T:8T8�V8(W2�b5dk|kHmDwm?~p7yr�y:V{5 }�<�@��,Ǒ@��8l�?$:N5SOXT0QXB�v*�~�~-�$� ${Q3�gz��NL�W=�h |kH[rQsS2u4�~*SO�[	g6q0yr&$`�Nm�NFOMO"SOo�Oo:P=�Q!�RL�R;So�Sl�Sa�SmT`T_�VeW9�XPY_eY6f[e�[X�[w�[�[o�[�\q�^>�^L�_R�`$KbY�blOez�eU�e/	g//gqhdhyLk8l$�lg6rq�s:5ui;uQLuQ�wnzhwzz�zGV{mM|7�|]�Q*�[��^%�JɅva�l'�\8�mD�l��hЏfS�^��`�\2�E�R�b��lfN�N/bS!�[;�_:�g1QhAGr�t?T�<�4�E��H��:�n$ 
N'NINT:NQKNI�N8�NF&OM�O]EQ_RN)RZ�S7�SU�SZXTU�T@�WR�WH�X;�YT�[$1\Q@\)^Y _?;`.s`]aN?b@@bH�b/te7�eL/fHnfH	gT(g;�hV�lLKmUwmP�rI�sLuB\uK�v-xRI{J�{=�~J�~P�~G�~2W�H��IKĉ<D���I�/2�=F�\b��B�TE�\K�V$FO5UO#lQ,bS5Y.*Y>�[,b;Ng5�~;~�3w�-ދ#� �l�-� 1 82 ;3 Y4 _5 [6 W7 \8 U9 VD Z$8 N?Nf	NZ
NFNKNJNPN`N0ND$NU%Nd-N1:NZ;N[>NdLNRRNe]Nb�N]�Nf�NO�Ne�NY�N8�NQ�Nc�N8�N>�N`�NO�NUOa
O,O`OCOOeSOTO_�OH�OQ�O?�OJ�Of?QaIQcKQPeQYhQ>kQ\lQRmQ]qQTsQBvQCwQg�Q*�QC�Q>�QW�Qe�Q[�Qi�QZ�QV�Q^�QYRP)RQ6RKJRdMRL�Rh�R=�Rc�R^�R[SRSYS_SA:Sf;STAS\JS_NSAOSTWS?bSXkSUpSSsSX�Sl�SL�SW�SQ�SX�SK�S?�S1�Sa�S`�SX�SZ�S;�SOT"TY	T]TSTO8TY�TE�TZ�TaFUX�Uc�V`�V%WQZW[fWd�Wl�WV�WZ�We�WPTXg^XP�XY�X_�XU�X[YEYXYEYN'YF)YW*YReYKsYZ�YV�Y`�Yg_[c�[B�[\�[a�[C�[_�[j�[>�[^�[c\f
\f\[\a<\\e\[q\Y�]J�]h�]@^Y^W.^Ts^Lt^_^N�^_�^[�^< _I_]:_eS_Jy_q�_N�_U�_e;`\b`W�`\b[bKbJ@bVSbHgbQibVkbevbbybebc�bU�bm�bV�b\�ba�bh�bDMcewci�cg�cW�cZ�cE�cR�c`id^�dk/ea9e;;ei?e)YeGpe[teZ�e?�e^�e8�eQ�eEfZnfbzfb�fX gQ	gOgbgI*gE,g@:gXag^�gf�gc�gg�gY�gN!hT8hF<ha�hlih'k5dkDfkZ{kR�kglOl^4lNIla_l[}lX�lX�le�l`�lZ�lL�l?�l[me%mawm6�mU�ma�mWn`/nZDno�on�oJ�obdqe1raireyrd�rZ�sC�sQ^t^uP0ub3uc5uJ7u^}vd�vj�v[�vJ�wR�wO�wJ�wYxTnx\>yG�yU�y:�y]�y\�ycze3z]zzR�zV�zc,{K~{c�{d�|c"}I�~Z�~a�~]�~:�~b�~&�~\�~a�~]�~R�~9Y	m`lW\�C�[�[L�aT�4��_��E�P�Z*�H~�aςU�\��S�Y=�fa�e��_h�c��e�A��T��b��R��9��e�C��W�V�c"�W'�b/�g8�D:�`D�W^�ap�b��d��Qƍo�lh�io�d{�e}�j��e��N��^��eǏ?ȏlЏZяNُ*ۏJ܏f	�d�T �eO�mW�im�cu�k��Y��P��f�dR�fǑZ̑^ΑSёK��^��d��]2�J?�<Ŗ]ƖcR�Z^�Ab�`�O��W��`ޘcߘe��Cl�NؚE&�oĞZΞaў[�[�D(�SB�bC�>F�]M�^N�IQ�TS�a�N*:N&�N6�S;T7(W,Y3�[0\3E\2^\3�]$^;�^*/f,	g>m*h�%��3Ǒ3b�7yr_!�O3�Q�[c�kKQ^#nf"Qh>W �e $�S7u!�v{�OSt�R�cKQ�R.�S�T<^X#\�_/g3�hs|"}%�~�/p�A؞5� T$!aNWSG�VUU\Y^�^L�v>�wX�{5Џ$ʐGG�ƖUՖRT{Q9h:u?����$6�N;yQFT>�V&\6B\�^6,gl6cw@x>yG�F�Fё΀ׂ�y(��e��	T+Y̑2��Q&\�b�e fm�~%�,��e�$)
NKKN?�NO�N@�Q�RNkS2�SFFURY"�[X�eIHhO�l9�v2�zP�~'jB�L9�U��P��J�l��SO�~�N)<PIQ(uQ6�RE^. _;c:�c7�eC>m)�m*�.�;ۏ'P[$�c�k%t
;uSO<lQ@uQP[F�e.ogH�Q=N>NaN!f[&$!T+f[,�c/f�y��%m�>�Lr �N(W�X.Y&tn3��=�Sb�NsQtQ#6R6pS5�S'T5�e6Bg1�m:L�ς6��B�N,FU4Zc[6e)�s7�|��>W�9��41 X2 W8 cV p� R$% N:
NXNMNeNANaNi"Ni$NJ-NR:N`;NZ>NN]Nm_NEpNR�Nc�Nk�N�NC�NH�Nk�N_�NU�NO�N_�Ni�NgO?ODOuNOeOOl\O]�Oe�Ok�OV�OW�ORPT:PFZP[?QgHQ)MQleQjhQbkQ_lQEqQYtQawQj�Q]�Qa�QQ�Q^�QDRU
RZRgRZ)Ri6RX�RQ�RC�RT�RY�Rh;SSASZZS^kS\tS\�SJ�SU�S@�SJ�Sa�SU�SS�SM�S<�Sa�Sb�Sg�Sb�Sk�S[�SjTPTIT2THTY4Tk8TiFTd�TH�TIFU8Vm�VL�Vh�Ve#Wt(WQ�Wm�WW�WP�W_�Xb�XeYS'Y9GYjbYmeYosY\}YU�Y`�Z=�ZpX[`f[>�[f�[Y�[Z�[C�[Y�[c�[G�[Y\Z\g\c$\n1\ME\bU\R�]F�]c�]_�]F^8^m&^T8^e�^c�^K_2:_\R_[S_]i_gq_d�_k�_Q�_g�_j`k;`ZP`hv`K�`i�`Y�`rbMbTbd@b]Kb]MbgSbLgbX~bdbV�bC�bd�b=�bY�bu�bU�bfcoPc]bca�cW�cY�cY�cKdWDdb�dk�dj9eg;ec?eOHe\Le\YeMpe_tee�eM�eG�ef�eD�eW�eV�e[/fMnfbzf:�fy�fb gG	g:gcgVg\*gf:gRBgjCg\Ngi~gg�gh�gj�gk�gPhc7hm�hg!jjck]gkv�kSl\4lYGl2}lP�l_�lb�l_�lW=mn>mMAmRwma�mZ�mZ�mknf8nEoV\om[rTurfyr^�rt�re�sZ�sWtVvtpuG(uM3u\7uhEuoYuI�ui{vg�v�vd�vT�vIwU�wN�wl�wZ�waxRnxm>ya�yf�yj�yH�y\zzU�zt�z^�zh�z`,{cy{Z~{e�{[{|^�|]�~i�~j�~m�~^�~3�~]�~d�~hQ<�_�_�RL�bX�_��^��_�_�k�c*�R9�co�az�^��i��w��c6�lo�g��Q�p�t=�jW�I,�j�v��gW�g��W��[��jƉi��mf�d��c��V��_��U��c��Q��D��O��^ċg��i��W�]�u"�`'�d-�J5�g7�@8�+D�4`�ip�\��Z��bэ`�X"�Pf�gl�Un�Uo�V��g��W��bǏ^ЏIя^ԏcُYۏ5ޏa	�N�V �hm�g�k��j��U��e��RR�fǑYёP��i��g��O �Q�i��l �\^�^�b�`v�d��mΘ]ޘ\ߘer�u��f{�WؚEў_�f�[�i�X�`$�c(�Z*�p0�g@�WE�_Q�eR� NA*N$MO<[O:\O@ZP7CQ<ZQ.uQ8T:�T>�V-Y<�YQ�YF�Z7�[F�[$\/B\8t^@b9pe�e0vfA!k l2yrYtHwJwD�y0�{Ds|7��1��DёG�Dy�:��A�5�A�Cno&��$6 N[NXNPNTN/NR-N-4Ne:NR;NB>N[KN[_NeqNi�NU�Ni�N[�Ne�NPO<O4O"O\PmZQ.hQMlQ:tQ[uQAxQ=�Q[�Q^�QjRjMRggR_oRT�R:SeASgNS^OS^ZSh�S@�Se�SU�S\�SQ�SO�Sa�SbTPT^|TJ�TCUbFU]�Vc�VQ(WGZW_�W-�W>Y8'YO+YPVY;}YJ�Y[�YY�Yif[�[@�[m�[X�[`�[c�[^�[9�[f�[\�[d\^\H\R1\a@\ON\oU\d�\a�]\^F^N^bE^K�^V�_j;`KR`c?adbSbWb[?bf@bggb^ybQ�b_�b`ch�cR/eX?e^�e[�e[/f_	gN*gmOgXhgfHh_�hV�i[1jlekcfkdlF_lB�lUmRAm[�q?GrALrQ�sbtX0uP5ub}vY~v;�v@�vb�w`,{bI{UV{ks|G�|k�|i�~>�~k�~h�~mbIT�R��^�Zz�h��n�^�V��b܃h'�lq�e��[W�Y�:��XĉD��Y��d��c׋f4�mF�Aa�\"�`[�A�c�e��fЏLޏB	�)�SS�^��K�,��JR�Cq�kϑ@��V�T��M�jF�Ɩ\R�_b�Ii�I�V��P�Vm�D�1�d$�f-�aA�dB�bK�aM�kV�nN9;N�NLSO<O7CQ.RL)RPWSKTETD�VHX8)Y?�YQ�[8�[:q\Hs^Ct^OMb3idK�e�eHl"%m�m-6q�s;�v7zz,~�=��LڋBl�:E�B�O&�S,�S3'Y5*Y2s^
�g Vn:zz3� �>�N�Y�YƉ3A� N�N,�Sf[2�c=�{B%�1*�#�5
N&$N*�S��8p�5N:�Q#�S�V4Lr5p�1ё'�{^�w��KQ
.s	B��e
ۏz�~'N+\p�$f[Lr�[�ONS-NO/OKKQApQEOSK�W`^XM�Y\>\GXbUTdO�e?QgS�g<hQtY3uF�vDj�S��1Џ�E�ƖW�9NNN\-NS;NS>NIRNLfNc�N.OJ\OIlQ`uQI�QU�QN�RU�Rd;SQUS7�SK�S<�S\FUd�VI�Vf�W6�XL'YK2ZMZ]P[f[Li[5�[Q�[c\Y\0L\Z�]T^Pr^Uq_U�_`'`-;`aKbN�bd�bi�c�cdDdRidhYeX�e_fXf@�f6pg^�gf�gI�hX�h=!j\LkN�lY�lS8nToGyr^�s.t[uE;uQYuP�vT�yK�zN�{V�{QGL�Hz�Q��W݄i��`ňAf�X��`��G��a׋^��f�]ЏA	�*ΐX�[��f�R�Q��OޘRؚTN�c$	�vNO,6R![r{|!�|j�($!N=fN>�N?�N<�P/?Q=�Q;�SJT?{TO�X	Y3}Y.�[M\9bBKb�e<�kE{D�A�Jr�A��"N7�N)UO�[?g-�gdkkp:�p5�~A��2�NE�NT�NUsYtZBz[W|^;�yQT��YVy'sYT�$�S/OS	�U�YP[�~P[ �N3�e9Vy(�~�Y�YZ l	7r�NM�Q3XT Xb8>mN�q��$z�� ?$�Q/�[=\#�^>�^0�eg3�zB��$Z�~'pQP[��  � FZ�N.MR)ZS/�Y�[/�^ K`/<y�~!?QHY!�[*|^w�N(SO �Y �ulQHS'l"�v�zP[���N?Q�Y��$�S4Y'7h+;u�v%8�(WXb"	g+h4>k(;m1��;7�6�R%4T%P[l(��-4�9��	-N �Rq\��Q��Θ?Q
�k �z$.NONKNI`NfNM�N;MO80RBMRH�RSTT/TWXTBXG'Y0P[1�[Y8^V�^VbCYeEpeO�eMgY/g$!h'9hY�lY>mG�pIuLuJ�v9�wMx8>yJ�yH�|M�~CQT�T�#��P��G��M��FǏQ��Ib�8��8��K��O?�YKN6P[ S ${Q.Y�laNTE�[00uF*� �Q�\#�b#�ly)��)�1 E2 B4 [� L$' NKN]
NVNONM$N\6Na:NQ;NBKNU_NZ�NQ�NW�Ng�NG�Nb�N]�N_�NdOdOT`OU�O8ZPa�P]HQQhQ$lQ[�Q_�Q[)RL7RgMR]gRToR`�RL�RZ�RhSTNS^�STTLTWhT`�TC�TDJUT�Va�VQ(WK�W\'YT*Y_4Yc}YM�Yaf[]�[W�[L�[\�[V�[X�[H\T\X1\T@\B^]&^Vt^]^_�_X�_g�_=�_L`d`g;`\R`g�`lb[@b]Mb`SbU�bf:cgwcd�cJgdg�eQ/fG�fb gS	gV4ggNgcag`eg\hc�kKlX8lN�lT�pd6qH1rV[rU�r[�sV�sRt<t3uT�v0�vSwS,{YI{Ls|a�~g�~b�~_Q`T�K܀V��U��b�t��\��U��a�QD�]b�P��e��9ߍ\"�M��Z��SُGۏO<�k��T��>�L��WёO��_�2�XƖ]R�`��c��Y��d��gؚS(�\5�RK�R�N,�Nr^�^/cg �hQ�U)bte5܀B$�T/�V/(W3sY@[bD�mD��;Ye 3u3�NJ�PAuQ.TOXT:W/�ZT�^O�eQ*:N-�N&�ND�N6O0GP-�QB6R+T/f[=\6E\�_,g%�p)��6+�-�3�)��8~�@tQf$ N?_NB�NIkSKTHJU=fUG�VE(W5'Y,\FU\4�\-cE�eD/f>chRm9AmJ�q8yrH�s4�s1�v.�w2�~_�Ch�B�25�,�;��Dl�(�.)�RM�EN-CNU`N@SOC�R1�S^(WBf[Q^\LU_T�`R�e�eC(gS�s(u7(�J��5E���/�BB��Yir$Rybt,�1����$��+ �?�NFU�[A�^F7b!g@:g+AmE�n>'�Gf�1n�IЏ2JT+^b3lb8�y,�~1��J��Q�S(Y'uQ4?e@�l�z$>N�^ _#�k%op.r$@g�v`lk�!$
N�S%"k%(u&�v#n�)1 W2 ^3 f4 f5 h6 l7 p8 ^9 sA sB �C }D yE �G $ N;Nz	N]
NXNQNBNGNDN|Nt"N�$Nl%Nd'N}-N>0N�4Nx9N�:NE;N0>NRCNnEN~HNwINxKN:LN~MN�RNbYN�]Nu_NFqN�sN��Nv�N]�NT�NL�Ne�Nm�Nq�N��NR�N|�NJ�Nq�N��NH�Nu�Nk�NV�NY�NT�N{�NS�NK�N��Nk�Nd�NO^
O�O�OWOW&O�8Or<ONOoOOoSO1UOw\OQO\�O��On�O]�Ov�O�Oz�Ov�Ou�O��OM�ON�Ou�O|P�Pf!Pv:PX>PwGP�OP�ZPV\PiePkwP�P~�PZ�Px?QoAQbCQ>EQnHQYIQpKQlMQgQQ{ZQ[\Q�eQkhQ\kQ]lQ>mQvqQNsQFtQZuQ�vQhwQZ{Qq}Qz�QQ�Qc�QT�QO�Q��Qn�Q}�QR�Qk�Q}�Q��Qh�Q]�Q��Qe�Qz�QF�Q�RSRtRzRuR[RYR}RORz)RA0Re6RP:R�JRzMRYgRgoRG�Rt�Rg�R{�RF�R^�R]�Rh�R��R^�R��RuSYS�SfS|:St;SQASbCSzJSpOS_SS�UShVS�WSeZSS`SekSOpS{qSksSptSawSv�S��SZ�Sv�S`�S_�SO�S[�SL�Sf�Sj�SX�S9�S_�Sb�Sj�Sq�Sy�Sh�SW�Sn�SR�Sm�S]TSTU	T�TOT[TgTPTm&T�'Tu/Tw8Tf@T�HT�hT{|Tb}Tb�T��T#�T��T}�Tz.Uv/UtFUPJUk�U��U}�Uj�Vi�Vu�V_�V^�Vv�Vp�Vn�VM�VRWU(W6GWaZWd�Wb�W��Wf�W��WT�WQ^X��XT�X��XlY`Y�YrY�Y>YW'Y?)Yd*Yq.Yz1Yi4Y:YxIYtKY�VYa`YzeYPsYOvY}Yk�YV�Yg�Y��Yy�Y\ZwtZ��Zm�Z�X[ef[_�[r�[5�[c�[K�[f�[j�[R�[C�[X�[r�[f�[�[_�[j�[��[��[��[m�[X�[6�[j�[P\�\f\B
\c\f\e\g$\e1\M<\�=\Z@\`B\rE\fH\�U\da\�e\j�\�]�)]��]��]:�]n�]��]t�]D�]w^]^|^�^`&^V.^e8^eE^�r^Ts^]t^kv^a^R�^|�^��^��^C�^��^��^M�^�^��^��^? _C_�_\1_�:_TS_`U_�b_]i_{{_��_u�_g�_~�_d�_��_|�_f�_w�_S�_��_� `}`�`k%`e'`r;`SP`jb`[j`��`��`��`]�`��`��`��`ma�a]aj?amb�bZbtbHbY?bs@bHKbjMbYSbdgbcibakbvmb�vbWybL|b�~bybT�bH�bX�b��bx�bD�bq�b�b�b~�b}�b^�b~�bs�bt�bf�bx�bx�bm�b��bv�bo�bv�b^�bW�b��bu�bhcgcU	cfc~c�#c�/cm=cXMc�Pct_cobc{nc��c��cV�ch�cd�c��ct�c_�cW�c[�c@�c��cide:dvFd_Hd�Td�id}�dr�d��d} et/eR6eZ9eU;ek>ed?e<HesQecYe8^e|be�ce�fe�pehte]�eH�e��e��e�eK�ea�ee�eA�eW�ei�ec�e��e`�eifufWfb/fH>fynf\of�zft�fy�fq�f{�fX�f� gKg�	g4gcg�gr(gw*g\,gg:g5BgrCgL\g@agoegNogLpgdg��gq�gb�gJ�g��gp�g�hChwhl8h[9hY=h�Fh�ch`eh��hc�hl�h��h�hOiz-i��iv�i�!jy*j�Dj� kw"koLkeckJdk}ek�fkd{k��kv�k��k��kR�kx�k`�k��k��k�lDlT4lQ8lpBl|GlyIlsalzrl�}lk�l|�lv�l��ly�lf�lq�l��lC�lf%m�*m�;mz=m�>mYAmhKm]Qm�jmwmJ�m`�m��m��mk�m��m�nunun�!n|)ny4n�8n^nv�n|�n�ov\o��oqkpbmp�up�~pv�p��pZ�p~q�dq`gq|�q|rz1rwHrYLrzar�ir\ur�yrSzr��r{�r��rQ.s|�s��sB�sS�s��sg�s{tqtn�t�uhuR(uS0ug1ua2u|3uh5u@7uS;u{Yuc\ux�u��u��u��uz�u�Lvw{vj~vm�v�v}�v��vS�vV�va�vJwwwbcw}fwu�w��wX�wu�wV�wmxd4x{nxT�x��x��xs:yv<y~>yV^y}wy��yT�yx�y|�yg�ys�yp�y6�yW�yy�y]�ys�yt z{z>3zXvz�wz}zzc�z{�zV�zr�za�z~�zu�z�&{�,{[I{gV{�y{r~{Q�{W�{jM|�{|�|��|N�|u"}|'}b/}oA~d�~��~��~l�~1�~u�~��~j�~]�~��~d�~f�~G�~x�~0�~h�~��~Q�~q�~5�~W�~c�~^�~n	r�nn)�4h:hQejvn��h��h���s�b���W��L�]T�EX������������S�����x̀z��K��1�yP���E�i�s�x�t*�R9�}o�z�b~�j��S��n��k�~�u�v'��I��c�go�R��a%�|=�sW�xa����kĄ�섋�t,�����Ʌ�}�b���W����u@��e�[h�]p����c����`��Feĉ=Ɖrf�]��3��l��Q��l��s��z��]��e��n��Z��j��hċlՋd݋pދ�勃�^�g�������m�q4�pA��a�w�[!�g"�<#�v'�Y(�G)��+�_-�m.��/��4�}5��7�h8�]D�NK�`T�VV��Z�q[�^�y`��b�qd��p�aw�r��q��d��@ƍ�ߍy�q�g"�f����nl�`n�{o�k{�e����p�����b��e��aď|ŏoǏfȏzΏ}Џ\яYԏyُ^ۏB܏�ݏxޏiߏ��r��q �n�}�p	�]�f���L�� �Q.��G�wO��S�xW�yc��e�|m�eu�s�t�����d��U�W��?M�xǑM̑VΑtёSt�^��q��s��o��fܔ���J��� �r�k��G�����-2�E6�u;��?�zF�pP�cd�hw�i��u��mƖNǖ�ꖉ �VR�U^�e`�xb�Qi���vv�y�oz�|{����\��I��9�����������Θcޘ{ߘWn�qr����u��Dl�op��q��{�T��R��sؚLĞkў��T �p���i�r�I�e��!��$�`(�V-��3�|5�8�xA�dB�JC�\E�eF�[K�HM�ZN�5Q�SS�qNϑ��&^$<SONkSB�WQY''YD�[<�]=�bG�vA<yI�~P��I6�R�Ff�<R�=���Neg�!R\2\2gbGk�~6ς�$#�N9�N#wPGuQGFU3�V2(W>�X4�]<:_Mb8�e@	g(l�vC�-��@��*�:j�:SY� � l�\
t	1 Q7 ^$< NHNXNTN8N@$NK-N+9N_;N[LNG_NV�N8�N:�N?�N[�NE�NP�N:
OOY�O7�OL�O\KQNhQHlQSsQ]vQ7�QT�QT�QM�Q]�QX�QXRX)R>+RV6RYMRM�R@�R]SWSYS_SFNS4OS`WS6bSUkS_pSA�S_�SL�SW�SW�SW�S=�SH�SI�S5�Sd�S@�S^TR	T[TUhTV�TY�TX�TS�U[�V8WP(WMfWZ�WQ�WSTXP^XJ�X[�XKY'YL)YYeYR�Y^�Z[_[Z�[G�[G�[U<\P�]9^W�^N _YS_AW_b�_HP`Ub`^aVbW@bTKb;�bA�bGwcS�ceidY�eY�e]�eG�e1zfZ gX	gMg7*gU,gJegW�gM8hQ<h['k5dk,�k[�k[lQ4lY}l[�lP�lM�lA�lR%mYwm>/nY�oDdq`�rS�sT^tY�t`5uR}vX�vQ�wP�wK�w_�yb�yF�yVFz_wza�zZ,{RI{[�|["}U�~T�~W�~b�~LPW[jZ�/T�>��^��X��^ςF�L��_�P(�[a�_��U~�E�B��P݋6�F�_D�X^�W��D��_яTُ4ۏAёY��U��_2�^?�3^�7�G��/l�IؚQĞTΞS�^�LC�IN�P$\�vW�-|T'8^'~b9h"BleQB^1_F8n$o�vH�5�q\$i�	�^	@g,D�8��&eQD�Q[WEKb!�{$< N3N2N6%NB'N^-NT:N1;NJ>N4�N_�NR�N+�NV�N]�N_�NX�N3�N8
OVOWO4\OLOO�ON�OQ�OC�OZ�OOPX\PLAQNEQUHQ[hQ8lQQqQAsQStQTvQL�QG�Q:�Qa�QL�Q>RFRXR[)RH6REJRT�RL�R[�R(�RR�R<OSMUSQ�SC�S:�SE�ST�SPTVTRT<T+&Ta/TN8T]�TL�Vk�VU(WZW7�W]�WQ�XA�XP'Y61YYIYa�YN�YI�[L�[X�[9�[W�[.�[R
\]1\C=\;U\Ze\R^V.^B�^e�^1 _9_T:_Tb_P{_^�_K;`_b`Ej`Wb/ibFybbbM�b<�bT�b@�b[�bT	cA�c^�cX�c?�cC�c\:d]�dQ/eF6eW9eL>ePfe_te^�eV�eG�e[�eT/f=�fV�fA gV	g1g\,gPegB�g[9h?ckL�kN�kZ8lO�lb�l_>m0�mVnZu[(uD3u\�vk�vRxOnxS�yU�y93z_�zK�zT,{Z~{B'}_�~c�~F�~^�~X�~M�~V�~ �~W[�I�hT�D��U�P�F��]��?ĉ_��P��Jċ\Ջ^�\�S-�Yp�YŏaΏKЏ\ۏ)�^	�R�A�;c�eu�M�ZǑ5ʑb�^;�cF�YP�\��b��Z��XƖQ �Vb�G��<��=�S!�c3�U8�QC�XE�XF�PM�GN�BQ�MS�X%N^!�_:�+N�$@+NK�NGO9O&\OHON?Q=uQPgRH�RU�RCSCkSH�SGT7�TB�TMFU$�V?�W/�W*)YDsY7�YK�YF�Y.�Y3f[i[)�[R\^;�^:�^Y�bC�c<	gDg&�hNckIfkRlP.lF4l>}l@n@o?upKdqM�qG�rN+sJt<uP5uM7u;~v?�vH�~2�M��G�J
�FU��B׋O�'�J	�IG�,R�J��Lߘ@p�T��G�� �ND?QHQ1�QTsY4�YU\A�]%t^pe	g3�g9uI��B�<�PP[�zN'Y&X[;^\�e!	g*gfk5lG:A �7(�/Ջ:NvQ<\&ё-$< N5N)NFNNN-N5�NP�NH�NE
O6O0�P3qQBsQJvQH�QN�QM�Q>6RNJRU�R@SL;S@USR`S<�SG�S<�S3TLTE�VFWT(W8'YD�YC�[K�[D�[O\6�]:�]N�^?�^; _4�_T�_Ab`Pb=gbK�bc�cG�eG�eK/f	g"gF8hD'kKdk1fkJ}lS�lO>mNwmP�yN~{D�~N�~S�AT�N��7�R��1�:��C8�N��Jُ5ۏHc�S��U?�MP�S��T��El�J �P$�H(�7C�=�Y"\"i`&�e�e��,*� N5�R1�_/�_�e�{$EoR0�R�W@\'(u,�lN1�N0OO PKMRBl6q(Yu',{&̑?��3��.ؚ@�Sc	g���e $%-N,�NJO:�Q:S1�S0�S�T/FUC�V �V@@\)�^K _�s2:y&<yF�zKȉ �9D�K��-�NW'`#���)a\B� uQ
N9N:S�[#q\;�]3Qg<�g=8h8Lk44l�l wm7yrC�z;�8�!!�E��z sY�\a)�l+�n;u�wWS$Ow� �V�nq\6qgRё?e�z��E�'R�1U;�VU\Uc9o*�&f�+��(;�#N�NR�NO!$OV\O�OTZQ<uQG�Q) Sd�S3�SETWFU�wUz{P�~ez�.��N8�RD�IЏDA�S�S>m�KQ�N)lQ7�S#FU5�W'Y4Y!�[.U^3f ����"�V NO(ݍ��'N?N;:NF�N7�N[�N?\OLZPO\PLP_AQ[HQ=KQZlQQwQ<�Q8�QO�QCRLRWR4)RT6RA�RE�SU�ST�S1�SET5T3}TX�TT(W.�WS�W;�XSYG�[?�[C�[I�[@\81\;�^% _3b_4aXb yb>~bXbM�bE�bE�b:�cM�cD�cM�cT�cI�dV6eJEe;fH/f<nfV	gckFekS�lR>mH�mWuS1uH3u[�vL�wHxPnxB�z]T{S~{E/}>�~I�~��F��Kh�A��B��D��R��V��Jp�SÍV�V��Jȏ[ۏ5ޏA�I�M��XǑN��J&�Q3�Z8�VC�X9NKO KQ;�R.�W.\+^9�_B`P�b8�b8�e�g+mJyr>{v6wM&{:�A�Ξ<^��ag$H�SE:W �[W?e<lAAya݋OG�OR�+�N
O6&O0�O2R(9S9	T9�W0\*@\'�b,g$�l#�p8��'c�%��1̑��,��)���T\-�!g	9�$�PkQ2�_u"�D�*:SH`A�eJg J�%�[7b	�RTXё!�N �V�s*N<eQ"0R<T,�V4Y+	g9egǏ>ۏ>��+�4MO $/�R�N,�R-YE�]=8^?t^;
f?%f<(u3��4ĉ0��7�>R�?{�XT �N3sY@�e!og2�m�q7�~3�~#�~5��8����2�9� P$$�NKHQIRG�S4(WEGW)Y8�[YePfKgFl/[rW�v6I{(�Q��S�<w�Ib�F$$�N �N3�N;�N2O<�Q/�Q>�SCGW,s^>t^9�^";`D6e;�m@�n<u@(uG;u1�|-:K��;8�5{�ۏ9�F �It�/ �<��0 �:R�7��2NN/�O:�Q(R4T8�e2*g"�z?Q;��8��;-�܏A^�$~�7(��NX[�yq_?QsY%Ye��؞ NGN\N:N=INHpN\HQU�SNJT:W1'Y�]&�^\id\�d	�l(�n\5u7wW�yS��@ň\�*S�:�<%N�N"�Vl"�2 >3 H4 75 *6 D7 HD R� S$ NENVNONTNO$NO-N>4N]:NO;NQKN9_NQ�NA�NX�NM�NR�NR�NWO``OXsO:GP6HQZMQ]kQZmQUwQ]�QJ�Q_�QERW0ROMR*�RZSRASOGSMsS]�SJ�SO�SR�SOTFTMhTT�T>JUL�VG�V>(W?�XXYP'Y:)YU�YR�[S�[T�[X\P\S\H1\M�\\�]O8^T�^:�^a _MS_O�_X�_P�`TbbbJ�bf�bC�b%cU�cYDdYFdb>e?�eA�e2�e@�e.�eL/fJZfB�f^	gJg&egNog[chXehX"kU;m18n.oQ�pL0qRLr]yr0.s>�v/>y[?zC�zaI{@y{6�~N�~W�~Y�>�TT�;�N��6�Uh�L��K��Q8��J��M�>:�?p�XُSޏL�V��L��OR�=ёQ�4Y�]�V��TؚLĞ7�I-�a5�L:�[K�LQ�6�blq\ 1 J$NE-NAKNK�NU:PN�POEQU8RUSFwSP�SN�TE�XO�YRX[4@\G�^GbD@bG�b[/eL6e:�hZ�sE�v2�vNzz?�{B�|MrS"�Q&�YD�9d�S�,Ɩ2ĞX(�JNFNE%NM:N:�NQ�N;�N=OJ\OK�OCPT\PK�PREQ@qQ6RERJ)RP6RC�R$�R;OSH�SO�S8�SITET<&TR8TR(WZWI�XK'Y@�YJ�[R�[K�[+\E1\E=\.e\O.^R�^8 _PS_%`BbAbA�b>�bA	cJ�cT�cL:dH9eL>eM�fA	g9,gB9h6ckP(u,�vCnxN�y?�z?�~N�~T�~2�JT�K�K��KՋG�p�Q��QЏKۏ+�O�;u�B�Q��AǑ2b�T��FؚP�T8�JM�MN�AP[B\yr�~$O$�T,�V,1j,�y5c�,V�,'Y �TQX)_�ebkl#4l�~$��)d�h 9� D$ NCN>-N@KNA�NI`OIGP#�SJ�SITG'TDJU7U[SY[P1\EbIMbI�bP/f=	g?�kG�v"�I�I�PǏ/��D̑�C(�LK�A�b�CN)sO4YHY�[!�]5�e4f%�g�l,�mz�:��4��!�N	?eJW�N)8O&�[�~��Q�$H�N6RQ�RG�SM�V)b*	gJPg)ehH�zQ{��J��.��w�I �7��X��]v�[A�DNG*NQO@�QLR>)RH�R0�RTVSM�S�V<�Y_�Y\NU\U^9�^M�^T�_R�_Ob@>e fWnX�nRoQ��N��-��Z�5ǑG�W�F!�7A�TB�DJ�8�Q���Cg
[OH:PBsQE;SH�VB'Y<ZZAd[H�[?}^9�^;'`D�`E�`M�bETdYe-l7jm<6rE�rG7uE�v�y'�{/�MP�M��B�3"�5�M��H<�5R�H
NM�NHeQ7�S1T>zfA!n'(uC�y=*�Jw�ۏ�R	Tg)W%V� ̑$P[Sf$~v)z�)S�-�R�V#zfl!1 J2 MD M$ NFNZ:NK;NJ�N8�NB�NB�NUOD�O\�OX*PVHQHuQ:�QC�QHRB6R:oRL�RI�R:S4`SFbSF�SQTR4TFJTMhTT�T;(W3'Y"Y[:c[Y1\P _B:_74bYKb>c:DdP�eG�eQ�eP/fL gL	gDCgHNgJegNhgP�hV�kC�kMl1�p*�qX�s=u=;uV�v6lxH�yU�yQI{<�L�Xh�@��O��H��D��O�.*�Wu�VяM�R��XH�H$�U%�T3�M5�4B�?E�K�L�O�VKf7egL�N@-NBKNM�N8�N2�N\O6RBMRsSG)Y*�[;@\t^-�_LbB?eLYeH�eF�e*gH6q6�~0�O	�"{�Y�I�"�P
6R�(g�e �Rba�'Y�Y/�h6l/op'�s35uhy�{.�~2r�y�%v�/$
$ZSim	Ux!NB�N6�P/OS4�S9�T�VI[W"�W1U\8^Bf$|i>Gr�rI�x=�{QƉ��Dċ3��*b�'�^ dk�N�_eg ��/ԏ)uQZZ-b!6e�e)g(z?z+Ɩ}TF}YEG� �>N2qN?�S3�S$Y'Y+}Y*�[2�[?\*�_"	a?a7?aA�e.nf<	gAmAя4��%ؚ2N�'OS#^ �@IY Nm�ek)n�s�W�_8:g�l&u#5uf�=o�Ֆ8KQ�V9�V�X!\ �]a,�e5�k-�m5/}�~>��-l�9$
N,N+N;:N;�N<ZQ?6R>�S2TD�T$�V(W;Y>]G�^Bb>/f8ag5�l(�t>�vI�Dؚ7$RBT:�T2TXC`8�bI�e6t�v,�{?��?��7@�(��?ޏ7�:qNIHQ)�[5\6q-܀=%�C{�1 &O <$�X'Y:?ao9 �EO�?����N$WS8�S;(W)?b;c6n"�v%��/�$l�?pS=�h5��
�fNaN;�O0�b	gyr0�u%�9�^ HN7haN2�[!�`�y$�~$�9�[�NR*Qe �
N;-NFCNRaNRfNK�NE�NHODO:SO7�OE�OGGPTePP?QTlQ=�QD
RT�RY;SKOSHUSRkST�SH�S?�SWTR�T3FU6�VR�VA�VK�WN'Y%VYCsYR�YR�ZOf[*�[8�[L\O\SU\G�]C^=;`Da6b8?bTybQ�bH�bM�b5�bR?eAYe?peS�e;�eF�eKgL:gB�k,l=4lQ}lL�l+;mHnQ~pS�sK5u<�u8�v:yO>y8�y=�zT�zK�|Q�~A�~@�~K�~>QGb?�J�@��9z�P��I'�[��F��@ċ@[�<��QЏ@ޏI	�OёC��C �U�FƖSR�K^�K�U��P��MؚH�OA�=E�>N�B-��N8�N4�NFSOA�P\qQK�QQ�QE�QQ�Rf�RU�Rk�S[�SY�SRFU_�[c1\h�]�chpeA/fDvhm�hHt(u^�vNcw[�~S�~bJ��f��Rň^��][�jۏc�(ϑ@ �Y �eb�F��K$�``"`La+���N'�^��$Y $�[%��!�[ p`'`d�`6q{k6q	l�
EN �T*�	}Y4�]�u"}!�O��S�`�_ s X$NBN-NENV:NNKNL�NR\OO�OA�QX�Q9�Q$�Q%RPRZ6R<�RVCS^�S_�SJ�SN�SLTM�T$�T&�V7�YS�[K�[U@\V�]Vv^O�^T _U�_O `0a<+aVHaf@b>�b"�c\�cY�cS�d@9eXYe,�eE/fCnf]	g@ag^eg@lIyrH�rT�v�v8w^wS�wEx=nxS�y]�~8N�L�G�N��S��X��T��]��^D�\f�`ۏE	�4ǑT�UE�1�`�s� N �O.}Y-�]'nfl%�$�.gR�lZ�O(uP1ZP%)R1(W%Sb(���+�[wzIN"sT&�V,'Y�_)?a+2k+��Ƌl�N&IQ"tQ!0R�S#i`2�`+�gɉ&"�R�N:N*�NL�NG�R4�RQ�SOT�TF(W.^Ea,g>>mJ�y=�~3ۏ/�H�U<\ '`	$zf�O�[��_Ŗn�$�� $1gR�f
!hB��9$-NO:N�NM�N6�R"CSIXT*�T:GWaWY<1\@t^5�b7Dd\�eM�qP�zc�H�G�]��W��7~�_�=R�C_N+�N�Q)1\*Pc>/f,eg31r&�v��(%NY
�k�p N2N9-N7�NB�N;�NB�OFhQ3vQ%�Q=S4:S=pSD�SBTB�V%(W0Y4'Y8\9\:S_@�_:a?�e4/f2,g/�g:'k+/n8w1,{9�,�T�>�%�;��C�$5qND�N�O1xQIRK:S8�SHT0�V@:W,�e �eB:g%�kE�rMeu	�~)QA܀70�:%�>f�0�H�E:�L$,{!�~ +v�Y�[*\�~
ؚ�S�SYM|�N&�NO=)RNOSIP[8K\-�]X^@9e*of!f�4��>�N:�ND\O1!PNZP5lQKqQAsQ7wQC6RF`S2�S/�S'�SC(W2ZWGY1IY;�[A�[F\N^\8^=�^FgbIb7�bG�b@cA�c=�c3	g k?qNyrJ�rD�rD�yH�yH~{A�~@W;��G��B��?��J��9�:�)p�Dw�Hۏ;	�?Ǒ7 �2b�,�:N�JZSP[�b�$N@NR-N.:NATNL_N>�N,�ON�ODR;�RDOSHbSL�S<4TChTG�T9�VL(W6GWG1YLT[MY[1�[=\?�])�]? _5b1�d>:gNg4�gG�hC8nBXoK�s4t �v&�~<�~,B�K�5ׂQh�9�F[�4��C��Iѐ9��>̑9H�7ΘEl�<ĞH$%O!R6VS@�S2sY7b:/f!	g��KQ N=N<�N;�N2�N;�N7
O6GP�Q;�Q�T6�[@�]' _0�bC^c?eg8�k?kp1t$4x5�y4zzA�{ �3%�4b�= �1ў;P�O�<7�5TX�y �{�bYuN&�