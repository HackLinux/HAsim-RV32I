�u��>EŞI�42�[�ח^�GG��Ĕ$���#EU��Uz�2���Ez�c��}�I���6����z_;,�f���8����No!��k����ǔ�u�/���N6��&
�Uz����ǔ�(ȹ&v�.�����K������W\՗z�G� :�Y'�˫:�s%�w��M�J������b���b���jɤ����┉�O����:��ݿ�`�ȫƸ��;��&�_�v��<�Nc	��ڿ]'�����?Q� �vA��+�l}�|b�"��<n�dGF��1�{��y�*�9|���q �\7�#���yD���b���1���E7(&��;�@��J�d�����0�s����p��x�dII�#��|:�>�1���<:�/sd&�bt$�o��P)lq`�`��+�p�xD;Z09 ���a�R5������ĕ�Z�V7����Z�f|E��+*��Za����5�������a '�0'��͜w^h�<YO,�'�t"�Ŭ_C=f`������t��e}�$Y�����@�� DK�Q����7�pz16�s������"�@���b���*x�B��S��o��DB/�g�D�\^uL�r'�h:a�ƪF}yv�[�`#P�-��R9�:6W��Z�3:�����SA*��l+����<��g������C����o1�3dM��B!�=�G�7�������)�^"T�������oA����A޿�A��c�����`RCIoy��3�%=r��ȼ��������� YU�~S�u��?8{���t1'_M2��3�B��4<a�~���ب�u��`z��W�#d��-�F� ��b�A01�Fd��$�� ����׍L���s��?W��y���ԅ�;_)�1(z�J0,[�iT��F=2�r��93���m��F�h;�1��N�P�#�Ϋ���Q��='�w��N�����e���q���ԫ>�w��XZ4�x�.��CQ 7ɫ4M�����h�ES� ���p��~��)�~Z��b��*;�vE�@�y��?��'�y���J�mH>����C��S�t��|���;�$& �j�/w��û�Ҹ�*Ms� ne�l�=w�t�!C����56��y9�;�3�F�v$a�-���`PPs���@��
?}�3<�1�a�0c0�5g�������'/[�JVr�սp��bD�m���7R�{�fos�?xf�5@Lq|���1��&H�~2����^�H4y|�vPÇ��^�� Ru\� ����E?����Y��\R����]a�ѯ�؏�H?F�ꦽ�l��3��	�Nz�!Oc�Uט;*�����g����jo�&��c�W�� 
쮠�y6� �(eI��w�	�V<�b�J�<1��dϔ����ɣb�i�H��e���U��0,Pf�����b�I�����k�_K_����D�_v����o���/7�}�;d�-5��֋�����Ȉ��H{�w�滆V5�Bo��S�sݚ�����ci[]����,{ �<��p_�l�iǣt�s�w&��a["j���,7�n�{����Gx�@���ե�#���#���`G���K�{؃���fv)�fv0�e":t�=�Q}؃�����
ڃ�s2�=�Q��`�9y&{�����`�Uu�h�`�g�k�e���`�l��r�(��U�kU��Z�=X+�eE�Zd`{�֚<k�<�f�*f ������0e���H������Z�ۃ�b9�ܶ*֢���5��U�&��]�ub�����6,�� {����O	g�w}��=�]�<������b���?�޵�����l��
"������]�P�][5��0{�5�%{�oX$�����V{ף~��kko{�ֳڻ>�}�y{��h���G�o�q�b���殨�mA��}۹��lߖ�+��2Y��Ǜ�:�~|)�Q�����-~�N��C�V�1��T� v6��