J�GLL�L�����M�LM�NNOO OPPQPNQQ�FMMRRSS�TTUU�VVWW�UXXWYY�ZYVZZ�[[T[X\\R\]]S]��^^__����``^a�_a��a`b��ccbdee`ad�edc_ffbfgg�^geg��hhiijjhjkkikl@DmmlAnnoo4EppqqCo��plnqmr�>ssrtuu=<vvtwxx;:yywz{{98||z}~~76}���51�������|~��y{��vx��su������_ ^ ����������������������������������������sr����������y���w�����vu���t�����x����������|{���z�����~���}�������������������������������������������������������������������������������������������������������] ������������������������ � ������������� ���������������� ���������������������������������������������������-(�����5 ���� �����$���������������� � ������������������������ ������������� �������������� � �����������������5 ��������� �������������� �� ��		

	 �: ;   ��!!4 !""##�$%%&&$'(())'(**��)*++�%'�&$�,,��--'�..//-,00./110221�334344556678867199::� 2;;9<� ==>>??@@<ABB<@CCADEEFFGGBDAHHIIDJKKLLJMNNOOMPGFQQPR SSMOLKRTUURJQETVTDVIWWXXVYZZUXYZP  # [[\\ NS]]^^$ __``aa]\bbcc_a^[bc`deeffdghhiig>fe?dih:9@;Cg( ' =5667788jjkkWH5+llj8l**kZmmnooppqqJOnngiorssttuurvwwxxyyvz!{{||}}z~��qp��������������z}~��������� % �������������������o�) n�����& ! ����������������������������" ��������������������r����st����u�{���������|x����y�~���v����w���������ON��b[��^a��`c��>=��PQ��JL��df����������������%$�5��AC����YX��������������������������m�"�����������������������������������������������'����������������������#����������������������������W(�����������������������������0����,������7� ���������������
���������������������������������������������������������������������������������������������  ����� ���	���		
 ��
��
��� � � �   !""##$$%%!#� � $&''(("!))**++&%$$##""!!%� #$� *))!"((''&&++*,,--..� %�&-,(./001122*+/2�33 � 44556678899::;;<<==>>7?@@AABB?@<;CCDDA:� �CEFF� � E9GGEHIIJJKKHILLMM>=NNJOPPQQRROSTTUUORSHPOLUFGVVWWXXMT� KYYQ8V7XW8ZYJ[[\\]]ZN^^__[]65Z4SN?B``^abbccddaeffggbahheiiehcjj� � dgkkllbmjcnnmgjmkln#d'hoppqqrroqssttuurvwwxxyyutzz{{||}}v~v}~�wv���~��x��������������������������������!������)�����+���������������������������� �������i������f���������$��������y����|�������$����������o����p���������������%���{z�������t���������s�������������������������������������������u�������������������������������������������������������������������������������������������������������r����������������������������������������� ������������������������������������������������������������������^`��� �� �  ���_��\6��		/+

	0  !!""!##$$%%"$,%�#  !!##+

		#$$&�3&�''())(*++,,--..*,//0011-0#!12233244/+55365+6#/4$+77886�99::�:
9;;77<<:<);85;=>>??@@=>AA?BCC@?BDDBEEDA1FFGG.FA=HHG FI)7JJIKCDLLIJK@MMHM*KM(NNNOOEOL�PP'P�QQPQ�RRQR�SS�TUUVVWWTXYY�XY��ZZY[\\]]^^__``[abbcc[`adeeffgghhiijjdfkkllmmg]ji^_hg`mabnnoocpqq1pqrrssttuuvwwxxyyv�vyzz�%{{||�}|{~~ut}s����}�������������wv�r�����������������������TWW����T������W�����pT�x�������wwxx�������~uu%{{~�����������������������&�����������������������������������VV����������oo���n������{{��~���d\��u���\��\���������UU�������������������������������������������������������������������������������������������������w����x�  ���������������������������������������n������o��k����l����s���c������p���d�����q�������e��������_����h���i�����^����������������� X����Y���������� ��������Y�Z�B���������D������������������������������  �������		
	�
 
���S����R�� !!""## $%%&&''$&��(('%)) #**&*++�,--��,.//0011.2TW33245566774�8899�100//..13WT22376655447�9988�:;;<<==:;>>??45<6..@@=/2p@?AABBCCDD117D930BEEFFCF8GG>:GAE@5HHIIJJ6KLLMMNNOOPPKL�2MQRRSSKP/.QIRQTTUUJJVV7WXXYYZZ[[\\W�]]^^W\3X__``aa10Y`bbVVccddaPY\MeffZOe[gghhNhefgfiijjghkkllekjilaQmnncUmdooppTpmnonqqrropssttmsrqt,98-buu4uH^vvwwxxyy_yzz{{||u}�+}#zx~~}{ )|]vw��~�$����%�|���(��S�H������wv������������"��z����������������{��!������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������-����.���0�������  � ������		

�����
����  ����	!!�""!##�#$$�$$��%&&''((%)**%()'++)*,,&,+����-..//00-122-01/331244.34566778859::9:;;<==>>??@@AABB��<CDDEEFFGGHHIIJJ?> C�KKLL��MMNNOOPPQQRRSS"LTT��UUVV�VWW��XXYY�YY�WZZ�ZXZ�V��[[\\�\]]�]^^�^U^�\�_�[_L�_T�_`aa��`bccddbeffggehii��hblmffbjM�kkllAAjmnnlkmoppnmo�qqrr�rKr�sttuu�qstpou�sBstlkundd``opiiggqc65ae7h8v?JwwvxyyIHzzx{||GF}}{~ED��~;��C�����}��z|��wy������������w�NM������PO������RQ�����S��9������������j������������}������������������:��������~��������{���������z����|��������x�����y��A���@���v���=������������������������������������������������������������������� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��		� �

  !!"##$$%%&&''"(!))**(++,,--..//+011,/020.*)23
1�3144�455�6ha776�88<7998�6:;;<<==>>:?@@AABBCCDDEE55?;BA<=@?>FGG58FG7�FF6GED9AHHII<3JJC=KKJKDK8@LLHLMMIM=NOOPPQQRRSSNTUUVVWWTX>?YYXQY5ZZRVSZ[[W\]]:XPO\^__``\NUT^]a`abb_^ QccddYVeeffS2[fggNPhhcdiiXhi`.-jjkkllmmajmklUnneng_*ooppqqb(rrqporplmqkorjsttuuvvwwxxyyzzs{��{|'&|}~~��������}w~}x�~w�������� ���������v���v������������������������������������������������$#������������������y����%��|��{�������������������������������������������������������������������������������������������������������������������������u����������������"�����ts������������������z��������������������������������������������������������������������������������������������������������������������������������������������������������� 	 			����	 			����		�								�						�
							
	
									��				��				�											
					�		��																									�			�											 	 			!	!		 	"	"	!		"	�		�	�	
	�#	#	��#	#	$	$	%	%	�#	&	&	'	'	$	(	)	)	'	'	(	�(	&	�)	%	�#	���*	*	+	+	�,	��-	-	.	.	,	�/	/	�+	/	0	�/	0	*	0	0	�-	1	1	.	�1	2	2	3	3	�24	4	5	5	[6	7	7	8	8	9	9	6	7	:	:	;	;	<	<	8	=	6	9	>	>	?	?	=	:	�3	;	=	�@	A	A	B	B	C	C	@	A	D	D	E	E	B	D	F	F	G	G	E	�H	H	I	I	�I	J	J	�K	�J	K	H	L	L	M	M	N	N	I	N	O	O	J	P	K	O	P	B	N	M	C	E	O	G	P	9	F	@	>	?	�F	Q	Q	R	R	G	S	T	T	U	U	V	V	S	Q	S	V	W	W	R	X	��Y	Y	X	K	Y	Z	[	[	X	Y	\	\	Z	P	\	U	]	]	Z	\	W	^	��_	_	^	�`	`	_	[	`	a	b	b	c	c	^	_	d	d	a	`	e	e	d	]	e	f	g	g	h	h	a	d	f	i	f	e	i	T	i	8	T	<	g	;	j	j	k	k	<	>	l	l	m	m	?	n	o	o	p	p	q	q	n	r	s	s	t	t	u	u	v	v	p	o	w	w	r	x	y	y	z	z	{	{	|	|	}	}	~	~			�	�	�	�	�	�	�	�	�	�	w	n	�	�	x	w	�	�	�	�	w	�	�	�	�	�	�	�	�	�	�	q	p	p	o	o	n	n	q	s	r	r	w	w	o	p	v	v	u	u	t	t	s	�	�	�	�	�	�	�	�	�			~	~	}	}	|	|	{	{	z	z	y	y	x	x	�	�	n	w	�	�	�	�	w	w	�	�	�	�	�	�	�	�	�	�	�	@	�	�	�	�	�	�	�	�	l	�	M	L	�	�	�	�	C	��	�	�	�	�	y	���	v	�	�	�	�	�	�	u	�	t	�	�	q	�	�	w	�	�	�	�	��	m	��	�	�	�	�	�	k	�	�	�	�	�	�	�	�	g	c	�	�	�	�	��	�	b	�	h	�	�	�	��	�	�	�	�	�	��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	��	�	�	�	�	�	��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	w	�	�	r	�	�	s	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	n	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	!�	�	�	�	4	��	�	�	�	���	�	�	�	�	�	�	�	�	�	��	�	��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	 
 


�	
�	�	











	
	
�	�	







�	�	





















	



�	






�	







 





















�	 
 
!
!
�	�	"
"


�	 
 
#
#
"

�	#

�	
�	
 

�	
$
$
%
%
5	&
'
'
(
(
)
)
&
$
*
*
+
+
%
,
TW-
-
,
+
)
(
-
,
'
&
*
'
.
.
/
/
(
/
0
0
-
0
1
1
,
.
1
+
2
2
3
3
)
3
4
4
&
2
5
5
4
5
*
6
z	x	7
7
6
8
9
9
:
:
;
;
8
6
9
8
<
<
=
=
>
>
?
?
@
@
{	�	A
A
;
:
7
~	B
B
C
C
D
D
E
E
F
F
G
G
H
H
I
I
	J
K
K
L
L
M
M

�	J
I
J
K
H
G
L
N
}	|	O
O
N
P
Q
Q
R
R
S
S
P
N
R
Q
B
@
P
S
O
�T
T
U
U
V
V
W
W
X
X
Y
Y
�W
Z
Z
[
[
\
\
]
]
^
^
X
^
_
_
Y
`
a
a
b
b
c
c
d
d
V
U
`
e
`
T
e
f
g
g
h
h
i
i
j
j
k
k
f
V
k
j
W
l
m
m
n
n
o
o
l
p
q
q
r
r
s
s
p
t
u
u
v
v


w
w
t
x
v
u
q
q
x
w
y
y
p
p
t
s
z
z
t
M
F
E
y
z
{
{
u
r
{
|
}
}
~
~


h
g
|
B
}
}
C
?
~
~
@
n
�
�
x
y
�
�
o
�
�
�
�
�
�
�
�
f
�
�
�
�
|

�
�
�
�
i
d
�
�
�
�
�
�
�
d
Z
Z
�
�
>
>
D
D
�
�
�
�
�
�
}
�
�
�
�
�
~
�
�
�
�
�
�
=
�
�	�
�
�
�
�
�
�
�
�	�
�
n
�
�
�
�
o
�
�
�
l
<
A
�
�
�
�
�
m
�
�
�
�	�	]
\
�
�
c
b
�
�
�
�	�
�
�
�
�	a
�	�
�
�
�
�	�
�
�
�
[
�
�
�
�
�
�
�
�
�
�
�	�
�
��
�	��
�	`
e
�	�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
_
�	^
�	�
�
�
�
�
�
�
�
�
�
�	�	�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�	�	�
�
�
!
�
�
�
�
�
�
�
�
�
�
�
�
�	;
�
�
�
�
8
G
�
�
�
�
L
�
�
�
�
�
�
�
�
�
�
�
�
�
9
6
�
�
�
H
�
�
�
�
I
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
J
�
�
�
�
K
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
R
N
�
�
�
�
S
�
�
�
O
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
7
�
�
�
�
�
�
:
�
�
�
�
�
<
F
�
�
�
�
�
M
�
�
�
�
�
�
�
�
�
�
�
�
A
�
�
�
�
�
�	�	�	�
�	!
�	
�
�
�
�

�	�
�
�
�
�	�	�	�	�
�
�	�
�
�
�
�
�
�
�
 
�
�
�
�

�
�
�
�
�
�
�
�	


�
�
�
�
�
�
�
�
�
�
�

�
�


�
�



�
�
�
�


�
�

�
�
�
�

�
�


�
�
�
�
�
�


�
�
�
�
�
�
�
�
�	�
�
�
�
�
�
�
�
�
�
�	�	�
�
�	�
�
�
�
�
�
�	�	�
�
�
�
�	�	�	�	�
�	q	�	�
�
�
�	�	�
�
�
�
�
�
�
�
���
�
,	.	�
�
�
1	�
�
�
�
�
�
�	�	�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
  �
		

 �

		�
�
�
�
�	�	v	t	�	�	p	�	�	�	�	s	�	�	�	2	j	 !!""##$$%%&&'' ())**++,, '(-..//0011-2-13344556627882699::;;7<==)	(	<>??@@AA<�>BCCDD>,	B0=A34@?5D9:CB;).-*E+2EFGG87F"HHII#J%$KKJLMMJKIHNNLOPPQQRRSSTTUUVVORWWXXYYZZ[[\\]]^^__``aabbccddSeff&Me gghhii jkkllmmjnooppjmqqn�nq�lrrssmsttqt�uvvsruvwwxxtx�xonz�kxooppjjkk��yyzz�o{{||p|}}~~k�{i��������}���������������������������������~fe���������������������������������������������������������������������������������������������������������������������������������	�����������������
���������������������+����,�����!�����N������e���������f  ����  ���� �������������������  ��������������������������������������������������� ���� �����������Z	���	������������������������������������������������������gg��� ��  �		

 !!""##$$ %&&''(())%