g���"���L�R�7]��>9�|�A�f�ϛ⬃�Y��>�MN��l��(�lA��t���w�}��{>���h��}���}��ӽ��x���z`�׭p��h�
�./\��*���9p͇+�#p�1���<~��W<[�m�p���)p*�u�ٹز�N5��T�� ���T���5�h.��������J���1T��	���`�f�T��LkU�iH�8B��n="L.�?�s������X�K�̀.-��#(*tD��0�\����[���8_ő�ը�������8�˰��ы�I��U�'W�[BJ�\���Z.�t��1S3e�������k��Θ: !�_�Q|0�=�s��Z���q�=�:>sH�:���Y�3c���Cf%��$�+�*Bfn�sK�p�h�o��Q$��d0��ϑ��@�߂���RD�F��m�!m�k�	�4���ȱ�y���zR��f���L�n����r=���R�<h�ro}�i��9_�;W��.M��ryU:�E��H�1L�l{{�W�[u�
�z�+4�C�����|J��=)�O�{D�x8��ZBa6�S�4�K7�?�SPl�5DYP�vJ�m��T ��"?��,�/����S�[rV-�7?�9���� ����dl�2�$��x�!�z[�ڻ�..7*��2+$;�!3+�1�5�dgtH�:�����_���ゼ��r��j���F.�ʨ��s�Q�?l�Q��\��?}�1�й)!�I�Ցؖ���)��Ƕ�T@;��اTT�����n� ���DC�Bz����3�^��ԯT�K�_Y��W����e�0K�n/Qj��.���"�p `�%�*2��c�h�C��V�����O!t�>F:��@��K�J���	�p�G_����zg�#��4,t6wp��I�6�h�]�~n����ᯕ����Co��S��0�r{����ʪ0���Jc��s���s���>�ژnX��w�N�w.ة(!^8����>,��xֻ���i�@-'������?`F�(�)�ʍYZXa,J�lcQ�f�2e�1]`�(�	[RQ
P]25����@�䮑V�q6�6�;	���d�HyR�N��x��@/@�u�1��rc��e,��Y����2�{x�+��[�"����] ؕ�c'��ys>�%�a��}��8�����.���WY���#������&�A��A>�C�37!~�ۤP"~�I�/�EP�w�0@!v�0J�_���a�~���{0�g%�ζUX�g���]))���*WB�s{�?亥e0W#�Ĉ�C���Ϻ|eB�@�%MJ�2_���[\h%�.��C8��>�ts|��F���(��e����7�WK~��K0��a�~(ܛ��z:s /����O��Q�K�R��]���õ��`�Y)z+��A�?_�Ig��+��ǎ�����ؕ'lq4<�,v�����~���s/�8���|��NY�ҿtv�
O��ʯ�ǹ�K%�G$�x�H,���1��:e)4�V���Zh����A2���v�º|�0U��8_
%�P!��#X �F����I�3	z��I[�@n#�}+Uyo{^,,�,�#zY�:��X��ADV~%�A��f�LI��p�W�C��̛�ؖ��d/R-����l���a����T�s�C�NE5��A�҄K�B]������ƺO�N)�~�v�gL4�e�m�g"��Ň��%��Bv�M��K��p��΍+�|2�%�)����ó�3��%��Y��-���ặX�˦�#&U&&;t&UL�EL*��D��MLv�L�L�9��,�ܜ�$db�Kg�`�����f�n �I���n�I��?�CLn�fR�Ĥ��d�Τт�ęl��d���D&+LL��LVX0�d2�[3��$&-&&�t&-L�L�*,�Ob�jb�_g�j����k&����319�3Yg�䏓��(k&�IL^519�3yՂ�̙��ܒ�"��ML>ҙ�n�䋉Ĥ֚��IL�21�֙�e��7�I�̒�IL6��ҙl�`rg�5�mr"�v��:�v&�L &c��̗]|����x"����'+Ę��W@� ��z=�>�ѱ���d4�e%V�Q//�p�Г�j�^��&�{/�a8例�c���N��>�iA���}5U($����9�e3����S-����X�<��`�F �pu:�v\��ڗB���� ��˚�K!i�_���v�a|���8>�L�����8��Ut{���k�&���޲����&ڤ�_�j�	����ɷ�&���Kg�I"ՉV�ӂɥ�ٛ®]����VF=4M���ʂ����N0_L$g6gb�Lm������S<k�G���3]���7"������!�U<b��W��i?�j&��F-)&慪gS�����?F#*	�=*�1*��Hi�q�hdj�9]�d1l�VC�y6;���{�#[��	$��u|��i�:�3�ϳ�k~L��{��e�5E�#:�Q���C�ze�(�,���O�p�a|�>`��N��Ʀ�O�W�K�I��,z�
���bnH�<�z�|<��K��G�L���e3m$���-����c��������vs�[;)��b̚9a�gd(R^@��C�n��m�x(G�8Ŀb����WRB��������*m�1>�ۤ*
����~�[�n����V��h�B�є��ѝ��Һ�4ʙ���Ff1���^H�::����ƛ����r�ݗ�O>6΀�o�U��㴪i�_]��s�዇��:�����.h�+E2\�2���Yq�FI�N�y=C�:��*�Պ=�/�\�_�(��ֿ�Dԓ׊(�G�|��"�y�e#�E,vŜ{3��#6���=����ÿ���P�&w�ji�`t��J/9��G.Q�Rze�����&��I��NL�K�甖�?�y�d�G�U�i�>�ea���L�f��>.4��� � ی�x;�N��*�)z��+0��4V��b`�� ��`���)�@t��v��0X*Β��K��0����S������U �Vb���9ܹV_"�qRqڹ�=6Q�����ks=����(��NP<����\:6�X�)R�Ok�!N�޴(_�o��1��H�ĶP�����Si�,��.�թ�<�{��X!�n��t)��r�hq��!����`G2�iK&X��B�K%�W��&�3���6B�2pF��N�t�z<�J��W�%|ļJ�Ln�K)&+$�)��������?�Q���7A�3ױ������6��m��A�C+eǷj�mY_re�����+D�#�uD���Vl��;�0<
X����7�����ט.� ��Q��h02��
�]I���Y���*�m�1�Oy�撔�͟��%�*�˪�}h�8��<������ЙJ��i�"���l���F�d�T@�31�؈��7�j�1.� ؑx�r΄za
̖�_�V���h����7������k8?I�8i�c�荛�	g�#��b҉�a"y��"����'�]���R(J��\�"X7w�փݰ��L���&�*�ò��!?O7��:�T�P�y<���j���_`
�K����b��呟���v,����ezKĳ��i����Fz\=�M�=���|	MN>.�3�(���l�2��.�������i�i��2�ri_�'Q//��/�5[O)rq�Þj+{:�e^���oׅ�o��f�;(^���s���N�4?y[�3�u���o�$�o�'�?=���Ap�v=
�A��-��'K{~��2�+�wv�＄��&�v�i�Y�gk���Q$���+A?�aN����D�G�=Y�N�E���M�`��>Ny����Ȳl��$3�E�kBe�(��R]������@Q
>wqY�A�Uf�N!UX�"0|��xө��MH��V�f�&����T&����}�����\�q�փ�v��e�gK1L��J��T��gG��Rvz:���x֛n��gX�)�[�%Fm���+�iE����"�)��`�-�؅Iw��a.���$��+��&���\d7T�Ƙ=�bb�9��?/�~P�ż?�����H�Se�OS|�@պA���"p`�Q��_�������һ���l��)Y��?�].�����ۿO�����?f�^~3��la�>�ۿߝd��ࡧ��� n�o�s�6_� �͇��6c�"a&�07���=��b�΍�ٝ���}?�f�/��@ :y�[lu�l/�*`�<�\t6<䖢��#�ڥH{z�v} #�s�U|K$�X�Ën�"[A����GN��aW�f�s5�������`�[�N�����Q	��g!<�v�׽ԡ\Jϱy?N7l�*���9�����n�4o��!�j}�p>���<��j��E竼�Ϡx�<��Z����}�>����� n��ԏ���C�v��>#]T����_�G��U$���P�4��`�﷢=�Mu^�"G��hpx�E�
+������*.ʁ�nɣ��;7��V����e��87B�ܰ�ٱB�%E����k_+E~�7�� _�4����;�~�"m:��u���|/�R2��� :�U}M�T�r����4w�"7	H�F�-"�d�M|{g�{��:׫���$��_R� k�)�	Bnݎ��������) �<:a��)��?��#�(��w�qxv<P#�EW�%���׹�}(3be�)eV�~v06�A�Mـ�e���~jót'-Ն���*����ަR�
�C�a�� ���p��
a~���=X(��
im{������c�R������@7���`��I�|���}̠/�_��FO�}��F��T��N�����P��4����Li,��x��d�-�<�KO���"�����iDB���u<���.�5��
�c2�a�W��
��AMrι��%W��es���%JHi_��&�R�^�L���{�x��� Y��^�X��:�v6���*3���;�Ҧ	�H�"��f��{D
4~u�=��`��6�C.Q�2����ݝ�C2�ȰC4�Q>N��M'�C���j�Ȑ��s��e<Hv�޼�{O(V����,���,�-��H��6���3e8|�&���zp���m6�ʎ8�\�����fG�m<�sD��ƳJ���Ƈ�|� �f�f� �OF�0�N�F�'����
���:�k�z�����*�������h��!O�[c%�Hjw�k(���N_�-��&` �}( �%0sR|�D��r��N�(�)��Wy��4�}���G�>:U#��r�jh�x��X$��^���~�2 i I3Г��K�&ᛩ�$;�����t�����_\������-q$Z��'�B��U=5�M�#�B��p���%IW39 �CK�}{|Tյ�H8�&f4Q�FA5a��df�2�_/4��mc2����؜�9�������j���w�W��*��<$	 ��DkO��Rη����+��? s��g���{��^�c�b;IF�ײ 0u�+c푩}&����AL}��^����~�l�t9es�H�f���[��5�<��X�~ȿ4Sw9�^��đ=+����62��0cG�k0�@��י��v�L���ܩ�+��h�앻��f�˭������h���M`�p��Ґ�$����M���Wa+Ӱ��z��=����=�9�6\�w��q$�'�dq�a�'{"�Vg���n��G�b^_���^.2̛��E�Q$2���PA�5�֝k~jˌ��k�O��
��.�<�
]Z5�bw#)�0U�Ц>�Ü��G�8�b7�+�E�{�<�{V耋�k�zm	`F�
0;?�yTH��k�3E���Q�b�'(1~��)�V��EBC���h	�J�!HW�S�@����%����E#% c.�8��~#��Ev�>�.�����P?e���~p�=�Ǿc��2sY\y��g��:�$��#9��=R+ǎ�#������,T4��PD�B�V�6N��쾧5YeY��'8�*^e>T�KV���rV9�W�
U.IV�����@`R�M�I}�R̯D���H ʹ��~��)�b_�Ӗ���
]h����P�P�ƞ}���n`�}����f=�j�Qhd�u�e����}�l� t1[��� vJ�tY��+|�<I������,_��"��-~
|�n:R�+0�Ѝ�ݑ��PR����e<��a� ��E���g���Yd�z�@#��:��p�fGa'�����Zs�����ո��W|��kM��KRCs��� �9���� ��
����~ř��{�Y5z�!6��e�-v��N�_Z߭��Fz{��JŠ,=]0�Q���I={��pC�kFcEo���}��D���}