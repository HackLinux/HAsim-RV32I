aB0��\�m�@��4c��}��G*;���4��^#	�ګɍ$f�^����\�K��ç��;J�t�*m?��$j�3l'墠�8�b>K	m?:.�}��t�#�� �yQ�"��9An�%�x�Sۜ�CL+�ة/OZ��&J|P�))O�K�#��t�����+�L����JCt�����΀-�5�B���x~[�A�S7ro,R6��U��Qs�K�B�aBIw!���R�*9��c��6}L��|e�Fn�k�VBM� ڒy��D�s'J��q��6ɜ�yDXLf�4mz��	Ω�Vk˞qa9u���W�����c�3�0��jS '�Y�2�q�$���yX"T M-f	V�t���ihj�7h�:89����B�'�p<>TW�ƹ*dP,Ԃ��P��nm����Uv��4�^Bv:vs^ܸ�||�ᖭl����T��`U%&��t���A`r$e�N3�p�5(�2P�S�ua
��nd���5ʝ?[�y(]l�PD��0��`�]�9�ws�F4�ј(B���m��beG��1�4k`C���@l���~�1e(�jr��.Ε����`Xi�K�K�f���,�U��X�XkT�2�W�Я�i�`d|s���H~���E~�����g$d�r��ڛx}/��nw���$~?�+bL������>qg��mŴ/�h��⌴�H�.���`��p����]R�KB~;�y*M02]no���F�s�:�BFr�Œv���V+�gųQ��7�\�!�].l/+��7�����)KW�fՒ��a[�\7���s�Ô��	;�P���"�zu�֣�,?y�{0������OX"��\�%Z[�N��L`�&�L;��ٛ�|eQq����
��������;i3��<0^�H�p�I�����nd�^�r$	W�H9d��kgR�!*��k��&"DwL�G��w>DiF��k�5$"k�c��S7m�Qm�Io[��"*5.�%"�ܣGnߌ�n�Qv�Ž�a�����"�5?;pS��9�G��^���BxF�.\`.\bGu�L�X��>�`<&D�}��`=�ǀ��a<�Ƣ�{�Ȉv��������S�r\��r%��D0W&O<�z�t��	��[t� :!�¾G�[������:t���WV��c��K!��D�:m�(w]��:m�η]��w��Q=��]H���'0�=��?����V��n�6�!{#��{NUu�I}�����\4�	���|��W�א�Y���9ٙ
t-�A�!56r��@��L���fGos8��[��]������3ьY�?����UF1.���X�c�l�x��NЮ��(�idǊSO�3�kK�8A؋�ڵ.��l^�ۿ�Xo����5>����R+sWz�%��-Ot�#~_��{�4&5�WQ�JS���w�(=5��KT�<��J/����}��o�s�[>J\�"�Gw��|j�i8�C|(��xCR`�`��8�B�>�Gu�W�[ێ�`����q	���'�X%B"�-V����1W)��a�P�"��NE�k9��q̼"!��#�B.�{�)���o0�X��ۣ]��f:�0�NTdMĸLV,�iG_x'p}g�0W����q?e�FuU5j�I�7O���b��@�6�������g�3v.����l<�ó�Z!��}c�f۶e�m۶3+m�֗��R��m�6+m۶�>��}����N�{v���V�ɵ���֍6�>-j,�<u;I���z���g٨�'�4l�P!�e����&��X*ێ�t�Y�>���*ӂӢT�~_�H�����t�ش�1v����AW{������q�'^*,���|�
�0J�g�hfW���а���&��D1�$�Ζw�{6 u�h���ʶH�U�[��͔��S���r�����|�lR��w&o�@&�G�]ܛ}ד ��5�ӼW��ۺ��,�Ւ�X^C��x�IJeg�<�[%������Ҕ�j�j5��z_G/�Ι�]U��C��nR�zF�j�x�U�:K� K��P�tM��a��1Y�1���	��?pg�R���L�NP��"kQ&4�֔�� ��Ҟ@[����7�.����Y���<U��HAmA#~���X"s�?f�:SE�i�lt� [��!����{2���e� P=!jӠ��0v��OZԡ�+��"�:p�R�pN�Z���@�q�/V�e��������h��?�Kɲ�U��v��Ȕ&�A�����<4�[0m��;FO��_@�K.�$��ͮ~x�|�O�7�nV!T�y�'��=/i�!����^ ��oh�>=Z�q+���g��/W`��q��-�c᥍8�+������U�Z���t�|� �	G����H U4S�ҘR�1z�_�b?j���).�,�1��yË��`R�<���]�F���z �]'H�K�>ep�)���Y(�nXZ*��*�f���/�2���JP2���s�03����C�tc��K�ʧ��N�쀕�0(���Lϫ'��7�'�{_�tY�}��>�K�i'�Krspʁ���m{xd{��&� �h_���P�^��E:�����љw�t����e^U�ļ�GY%�Z���t\�i�YKXCn�f�~Z@ہ�P�lvB�/�L�JKC�}]�jp`�r(ޱ�Mݭ�{�]������yg�?υ��[�!ȟ�s�<�A�B�P���q�LH0��o�B��z�_�:��y|Z�q�����J�S��m�A�6�V:*��^*U�����=��j[d�x,������OM��$�;ڛ�Zx��9�XXLIE,����?8f��8��_�+���ʹ�j�" �d��f�F���X#�2��6�lֺ�,��.^w}o��ݏm,6ikX�y��3~�|�m�{��2=����ܺ���{|>���(��o��U�d��4��>��D	����Z�2EL��+��m7��U�"�)���y��%�(�<FrO�hT.M�֛��E3 6yͳx-�p:��ڜ$W�x$�׼f[X�D���[�5�k���V�'�_�z�/1��vh1`�`ٺ��V�_rh����A�ת
Es���Y���ex�ͷ݄�`i�b@������F�r��	z>d�"/�
��A���k<n���r� �IO�(1�0��J/��� F��1WiP�ީ��/�}(}�)��u�������xjd�`��T�Zo"��S��9��EGf�΋�l��h*�F��ӈ�zu0��PS��6���sD�/�G���XZ��UOp�+�ME�l9���D��$�ej)�j&�HƄV۾�����e���#e�IF�5'���J��"A���r{��|#-wt���RN�	����J��p0J:a����F|���ñIB�yT�Ru1�[I{���;�r��=�ٵ�/o$�M`
������hc���Y��s�>�	#�k�������F����)����F;�n��#L����#���_�����N?�1�`
C����%`�X��hy������u��w'�&i�����Xaa�Q��L��Z�I�er+�0��+�,�pO��͓����fe[�]��궵c-��pÔ�Q|[�X�����]|����pL�΂�Pa��FYb݆9���{�J�c�ø�I'Xg�����	�s(� ���v�.��t|E ��9V��y�j��������+����/�\��[��O��k�3L��d	�&F�V�f�X
wL�N~���z���2��ɮ�2��g�� G��ꑓ�B���qxA��IN.����O���� ?~hC�Sa�/�Q��ɿ�
ʧr(����AÂ�y����y0��4c�s��V���LC��E�X��iD|��P�a;8/�ݾ��` QT�G��Nݗ��?���z1� f�}��!�w��izq���32�g�˰҅q�b�PK��Y���-V��,�Iz��x�iW^ZT6M�C��
�TDY�L"R+�t��0U*�L�x���ʋSR�M�L��\��XL�ߣ�\Xu�Z�\e�c��Pl�M�v��dd�� h�M��&���^x�}�މ24��1RM���'!Oj�8�G������K�
���_�A��T������n���CkC�t����E C�ͥ�Q���Z������t�A�=]�+��2��k�Y��=�Q�²ŹxѺjx(=|�����M$��o�?n�_��o��虝�U�����NO�F�`���*b��A��m$9D�`=��1  ���!q�o�$3�JB�ݨ�A̶g�d�͖�j�Ăb����� �P���R�+�c���:������e�9!u^n�⁅�5i�zvEް� �u[a�~�P�00b��5��6Y�
pJ�2ϧl~1O��%4H�A��/o}��������#Z%�ۚ�MP羇�p;�tw'�.��ص��[dC�*�Ѷ