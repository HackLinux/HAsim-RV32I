��sMBv!�1f> e(������'U���7K��*~�ځ��f�q��_�}�~�аcu�{��E�
�?�rQ<-UJ�{�e�κzZr�k%��i?�˫�<�.�k~Z��,��c�V̠�Y4zН�O���J�A��� ���>��tE-�)�q�ϛ*�yM},��dm����JG�lr�]3<�Ƣ��שe��2L���_�&�%+Q���E(�T��t<o<VY��z��A��Jw�V�V��L/�������1�t��\��7�jU.�&��eV+-�@oOJ��M����$��e�S6ŨN�^�mu������d �$i��ީ>e���I4E�5�8xO��n9�b���~����ޠ�w�ꎌJ/W�<ݺ�`���_����X0;��[M�h}�V�{����?W�"�j����W����8�����EG�H���YCW��[����}9����I]l
��W	YA�:%�)�ʧLwAm~�=P�Ry��=��r!՗�V���%���I���=vR����ťH�q0j;�r������xM��b�Z���V+��+�g�ڞKuQ�,Е�fQ��ջ5��z��B��T�@bɾ�)	�B�uD�������a�|*���*��G��oN=�ҮS~�W^��&ʞ�n�=�i�n0,a�ݰx������U�3?�;]	Ey��b�f��NlA5��+s��M E�l_��g���褨֕T�H�ޟ���U����
B��m��4/[�`��(�"M��.��K��a�?`I���%���#n^Y�k!x����ҒC�;����,�V��T�ȷʼGj�N��R�zW_s��j[���������+�,$/VD���(b3�&����õܳV�VPPE��h��HsT�V�Z�^
�4�@�=�yS׮��dO�t��]%~J�mۢ��W�񳀜�ATo�Y�9��sFC4�*n�(NV��!��t��TGp\U�%u�To��)L���
�h�z�|��>����Ī�|!W��x���7�j(>d0��?��z=J ��8�� ��V�Ͷt�z��mY�l]6J�����=�o����֝`��f���y볂}H���������Y�Z�Qש�;
��y��uќ�z��Ƀ>�䉿�пL+~�F�?ѫ�Tt|�Z��tb^�w=V(�ת�������5�qiȳ<�7iU�q��J9wzBR��*�WT0~��1�`���Y�k�TݳeJ�	ah$���(�W���|6�:�Op����#�̿������q	��T�]=ش���k�l�=�2���RtoH��w��Eb��pg֋�k�E�N�ݡ<�� 84�gؼ^݈��q�Գ���ݎ) �q��#��i_��b��g��dl��,ɪMx�	Wf��):�7�rM��m�8Bq�CrC�%�)d�Q�'�Z��8rp��H�����(��9ҷ'�P�JFO
!&��x������%��6$�'�����+��Xd>%��p�]:G�ˢ�3t�69�(��	z�ǖv��y���sGxq82�Ċf��8�pywsb"�a='�7�ז��F��p�=3o.8�@�Ǡ��a�1�2�N�1M�L3S59 ���~Doq�Ť��#ia��ʰְ۱q$Jǜ�$s�s�e�_��^�<����Љȯ(r����a���c�a����dSv�Ŗ��1��=�~��>�^k��:�ǽ�R\y�}^~�|^�[K�#@��n.�.z��g�-):Fp6����m��ͻ��=#�=F<ٹ��u��O�+tz�/�c=&�d����׿i�tN̓�W��Y�r�v�ɚ��|&�4joo��'l���%^u)���GSC�tu�!c5aA����3�E��=ɪ?��ɽ�V!p�K2��#�[D��v��D������׽O�]�_��p��X�d)�))��L3��1nV��t[�M��ֆ�=φ���<��ɸ�.h���	7.�<��xE�Օ�7H��vy�F`Eo���g���z������[ hc�n$�qVܽ��3hc��:Ćxu�c���/䡎�5�w�̳M���2g��򲲍�o���VqKlu�]}�Dw`��p��5[K���U��+�����ް�P���r�MV���F��\��;�X�.��j��.n��K�K�K�Xf?���c�;�;�;�8��t�l����t�LAN`�d���>��]g=⵿���f�����4ş��У�f�9���������L���-�/3��Ƹ�ھ� �c��� �����[�����	���P]�B<�CM���Iؙ%�LY�E.΄�:�u��c���h����������`��Ѥ��������(�M�%&`���k���lϏ3��X�8Ϫ"�VA�D���HC�x�³L�T��2�h��w���{�3��&�2诊ZW������fY˕u[���.^V�ɟ�E������8٥D�D��#�Ǽ������٪a�B����LY���Ñ~r!���Vl�'Z��́� [o���#	�қ󵪝�91K��@r�`�����٩�U�gxe��}>n�>i6az��h־�[�UD���Zئa{�Ϭ;"w�qfѬv/IK�z��:Ǧ���d_�|1��Pد菀$ҨY�w�q��F?�͈��ꄼ���;n�Y+f��06�:��-�&Y��	�����Z:I�w�^�Yn�8���c ��&�L�3c��@m����Bw҅��(�N�W��;F\�<;�PNMߺ�� �l^]��i��:�o���c�Q����ԃ���1�����ި�$.qى�6�"��?�4@��ܛmc��:6V�0�Υ?7���(_U�cF�e�,��G����-Zg�+)����Su��gqq[�Jf��\睅���P��.��K��]���rl�	�����������w��,<	V�����I��oS��,��,Yr�z�o��)�;�	E��Ā\]D6I>�V-�c<Ն�{&E� !6�A��>��֛���f���V<<K����_�C����*oj
s��*3{��
�3Ɛ?���^s�28y�ƈ��-(�ٽR6���cm�6���-uc;�ͧ�bܰ��L����q�	ͦ-�f�"�g�,F�|�t:A{�;�/J��E�f\!vY�L}�����M���|۟���zS�S���2�M�)�Z���%.�;��,�0�% �s��<�}P��l��N�Ѣ�9��ˠۢۨ۰۶��������6��,��l�����&�$�����4��	�9�aX{D�R�T�\�\;�:��\n���c�c�c%�r���P�*�J�jhz^�v����:�q�s��f:�!�y�s⵲q�cs�����`�si��i��V6o���XF�ڜ������\��X]1"��3ȳɳ�o 626�.��͟��g�cO�Y{�����޴,j��?�o �O�ޔ�g��/d!�_�i3��f���f���c.+W3ה
&�1�73O&���/�!i$%�Nq��Ɍki�t�Л��d9ʂ��7�̝�q����Q�z�yov��g�M��ٛmhg/�ܽu��wM�~���=ǅ�k�D8J��u�s6\;�u)(��葍H]�B��50�'��Y�p:�ﯷ�ٖ��3cv,�m=����g2�o�q�;f�h" ���~j.�T���6e���`=Fc�q�Yev����g+�T����o���-���oV���2Ԟ���4��G�/�XX�c�"$$�Bc�2c�N�j�0�[L�Y�n�V���ΪA���amg��1���#|�l*|Y<��B}`��դ��������dƋ��Uj��Ǆ"�0��Rd�=I���r��*����;��v�G���{e�9��͢
_�J�!qѫ�P�Zz������౪�.��O���v�u�ǂ���qHJm���K�#?޶���X{�i��U�"<~c�TxX�J��$
�b��e?�.�Y)�Y����Q?`�}�+ؙ�@��ё�c�7��B���&Nm��p�x��Żww�BA|�V\J������Kˍ�׳��%⛭]5}�;w���l~�m��.Q