~r�|�|��D|�܃��� z	�WZ��^$1*fd�������i��{�G,i��O$��'��H�W��Y3����Z���'�z�y�5򞷭nf�]�����25��i���XT|'���$�ޏ���������8��rg%��PR=�^�[$���A7x�Yɤ�5���`v�˴<k�u�u6��8r�9��t���Aޮv��ݜcߌNz��]�=�#蒩�s΋�F����0�n����]�}�=�Ǡ1ڂT���0"E#m��Ri�<A�O��Q�Յ��崳��4�C#W����я�3���5��(Z�#��3̙�l��n�`Lj�J�x:'~�3�$'��38���{�}�]�J�J���N	�����|��!K���s��Sn=��mw���no/�;޳��~t����X�����=P�W{��.�go<R7���@4W.-Ai�D.׆;ᚨ�[O�KI�x�h�bxE��^�!?H��t$�(5t9��򉒢�.�^ćF�؞��s����tҌ۸�����_�g��_�J�@'؝�y!iF$�a��)|�Gp�Nx��P�Q���m��j��Ờ�{�WQ��RoɦE(���������,y����x�|�r�*����� G?w|3(p�a�#诶��Ţ��㋗���x��4db���B~�����H�
�V��M�z{�WLZ��JBC��V����\�H&�]Af3�ډ���pZ�$i���߳��/��d��Β��O�Ϭ)�,�g�Хo����ϑ��)�p=�%F=��s�z�X�>ͦ�h���@`ߵ�<�1&�e���Z�~�<,B�/"�x7���U�i�#|O�����AR@ͤE웘�
\Ƴ��7m�9mw=�[�s]�d�&�u���"���5��HsD6�-y�a��h��M�%W�G�7GZD:�I:G.�״g�=�@=�a|�)M�ᚤ���<�ҏ�OП�W�