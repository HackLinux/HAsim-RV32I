���^�^������x��Ԇ�B�B��چ�ϳ����ؘ�س����س�س�ز�����ѳѥҳ�����������������������x�������������x�^��<��@����F����A�������^�����Fx����FF���F^��^^�x�x�xF��x^�F���^F�]]z��ffiiiyyyyi��yyiiiihhhhyygk�m��nzzzk�����N��`�����!�~~~~~]~m~�ccwcs�~~~�~mmm~~mmmmm~nmX~~m~m~m~mm~~m~K\�wwcq~n~~]Z~~Q�!�˲���`�iil}���nzzzz~�̃��ghhyhhhyyyiyyi��i�f���aKZU�{t�   D�bP]]]]]]�s�ss�omX��������c��gyg��mmXo�onz�h�eee}uupiiiH[b�j����|���ӺӚ�C�������A��x�A����t��x����fauı��������e�����}�����{�{��}��������f������ܜ�_dd�w���x��^�^�������x�������L�����ѭ��ؘ�������ز��ز���ز������ј��������ҥ�����������������������x^߆�^F^���<F�F@�AA��<���F;FF�^��@��;F;�^��F�^�^F��L��F������^�^��]]U�����i�yyii���iiyyiehkhyyhlz�m�ݍkkkzkn��l����`������!!�~Z~Z~~Zm~�ccG�s]m~Y~mm~~m~mZmmmmmYZm~m~Zm~Z~~~m~~\�wwc�~~m~]~]~mQ�!;˲|������lknlz�nzkkn�҃_�}hdyhgkieiyyii���f����Z]Za�{�D�DDtRbaY]]]]]Ks�sssc\XVV��������gg�mm~o�~Zahie��ff�zrup[KPlHN���������|��^BB�^Fxx�L���������t�t�L��u��fn�ı��������e�{��r��������{���}�r���y��������ܒ�Xdd�w������^�^�^�x��൙���ʵ���������Ʋ�سֳ��س��س�ѲѲ�ѳ�ؘ������������������������������������F^��^���FFFF��������BBF���F���^A���;;��^�F���F���xF��AA^^^�<����]KP�N��iyyhHiii�iiihyylkkkl�hzn�o��nkkz�nn�ll��N��������!!�YmZ~~q~n~��cw��\~~Y~~~~mm~~mmnmm~nmZmm~mmmmnm~n~mY\�wwc��~nZ~~qmmQ�7�||�`���l}nn��Ozkkk���cgnnlll�kkhyyyHii�ii�����Z]ZU[|RJJ�J�{baY]]]]]]Ks��u�c\\�����~��g_�mm����y�f�e���h�Zruu�i]SH[�����������˙�ʙ��Et�?��E��x����E��t��酯�fZ�ı�������fe�������������b��������iy����ī��ܒ�_dd�G���F��^�^�����xx����ʵ���˺��������������س�γززѲ����ј������������������������E��������������^߆^@F;�<�@����A��x������^;��^�xA���F����^F����x�x@��@�AF��<��<<;]]q��ii�iiy�i�iN��yyhllSg�kzknmn\��ngknkkn�}zl�����`����!!�YZ~Z~~~m~��cwcs\Y~~~~~~~~mmnm~���nmmmmmmmm~mmn~��wwc�~mZ~~~ZmP�!˓������lzn~��nknkk}˄nmn�kzklgllhhy��Ni�iN���ZKaa}b`j�j�j�[aZ]]]]]]]Y]�\�s��\��oo�mmmm�gy����yyylZ]]]KKuu�p�inHePuu������{�|�xLLxLA��x��x�x��A�E��t�x�b�f~�ܒ��������i�����������u�������u������������ܓ~h�d�GԵ���L��^�������x��������t�����������������������Ѳ��ز�Ѳ�������������޹������������t�����E����x��<^���xxx�xx������^FF�^���^FF���B��^�^����xx�xx�FF�xF�������]]Q}i��yyi�y�y�iy�ylyhlhhSk��nmm�ҼnkknnOn�znll��b������!7�Z~Z~Z~Zm~��cw�s�~m~~~~~~mmnmmnm~~~mnmmmmm�m~mm~\swwc�mZ~Zq~Y~u�*���|����llznY��Onn�kkz�~mmn�kkSSllylyyy�iy�����Q]aU}��������lza]K]K]K]]KK]KK]\\YooXm�gdghggkZZ]]KK\K]K]]uu��}�NKIHU�������������x��xxx�����A�Fx����E����x���fearĽ�������f�����������������������������ױ��Ċ�d�_w�������߆^�^��������L��ʵ�����ز����������������γѲ���������������ټ�������������������t��������x^�^^Է���x���AL�����F�B^�F����xxF������^^^F^F�F�xx���Fx��^��<���]]Q}�iyiy�y�yiy��yhhhllghgk��nmn�ـkgknnnn�pZ}zl}�������!�QZZ~Z~~m~��cwcs\o~m~~~~~mmmmm~n~nm~mmmmnmmmm�m~�swwc��m~ZZ~~ZZ��7Ѳ���b�}zzn~�znnnkkgn�v�nmn�kkghhlhyh�y��yiyi��q]a}}llll��lll}zZZZZZZZZZZZZZZZZZ~~mm_nnnnZZYZYZZZZZZZZYuuuzllyihHHHNii�W����������B^^^<�����^��x�E����Lx �pedku������������|����������ƭ�������Ē�����ױ��Ās�dd�Gx���x�߆�����x������x��ʙ����ز���ؘ�������ֳ�������������������������������������������������xB�^����x������A���^^FF��^�^�FA��x�FF����F�^Fx�x�xF;�F�A��^<�^��]]Q}iiiiiyyyiiiyyiyyhyhhgkkk�nnns�kkn�nnn}}Zazz}���`��!7�Q~~Z~~ZZq�scww�~~~mmmm~m~mm~~mm~mmZmmZm~~m~n�mm��ww�qqZZ~Z~Z~�77�������}zznq�Znnnn�k~��V�n��kkShgyhy�yiyiiii�i�Ullll��l}��l���ll���l�l����l��ll���nnnnnzanaaaaZaaaUaqu�Phyl��gdhh�ly�f����������Ӛ���C�F��F�����tt�x �zedH�ƽ����������ı������������������������ı��ıreg�\w��Է�x^����^����F��E��ﵵ�t�Ϥ�������������ֳΤ��μؼ�����������������B����
������������t����x^���x�����������A��^^������^���F^�^���^^���^���������xF@�<�;FF]]Q}iiiyiiiiiyiiyHyyyelhShkk��kouՍnknnnnm��~Zz}���p�!!�QZ~~Z~~m~�scw�s�mm~mmnm~mmm~~mmnmOm~mYYn~mmm�m~�swwc~~~Z~qmQ�7!�[�}}}zZZ�~On�nnkm���k�n�kSghSyiyyyyiyiiyii�U}}}l���l���yl����l��lllll�ll��h��zZZZZZZZZZQZZqYQ]QY]qu�qhhhh�g��gghhyi���jj���������CC�^^�������������x��qhde����������������ı��������|�����������ı������legdw�����xÆ����^���������D����������ز��ز����س�ҥ�ֳ�����������������Ȇ����������������������x^�<<���   �xL��A����FFFFF��F��xA����߆^��^F��FF���^F��F��<�FF]]Q}yiyii�i�iiii�eyyyyyhhhkkkkkV�J��k�nnnnz�ZZ~�z�zZ�!7�qZ~Z~ZZm~�ccwcs~~~~~mmm~~m~m�m~mmnmm~~~~~mZmmm~�swwc�m~Z~~qZZ�!!�naZ~ZZ��nnknk�m��cnkk�klhhhyyyyHe�iiyii���}}}}}}}}ll�}���ll�l�}���lly�h��lha\K]]KK\KK]KKKK]K]\Qv�qhdhhhhg���g��yi����������CԆB^�F������������������˄�He������������������ǳ�����������������ı����פsfeg�G�����L���Ԇ�����x�����t����t���ֹ����������ز�ֳ�س��ֳΘ����������Υ��������������������������������x^߆����   D�x���AF^^����F�x�^�xx����^�^����F��^���x�FF���^�FFF]]q}iiyy�iiiyy�i�i�yyyyyhllzkk����a�nnnnnnz}~ZZ~ZZZa~�!!�u~~~Z~QZ~��cw�s�~mmommmm~~mm~mmmmmmZm~mm~~mm�mm~~�swwc�~Z~ZZZ~mY�!!�~~~Z~Z~ZZlZnnnnnnm|�wzkkklhhyyyy���iiiyyii�Qa�}}[���ll�l��zl�llll}llll�ll�ll�zZZQ]ap}paPqaaaaZQrv�r�y�yhhh����l�hhy��������B�Ԇ���������������������E�Յ[de����i�����ī����JJĩ��ؘ�|������������������r�fd�sG�L�����Ȇ�����÷xxx�����������������������س�ز��γؘ������������������������������� ������������x�������  E��8�x����F��^��FF���xF�FF^�����^F�x@����F��x�FFF�<��F]]]}���iiieiiiiiie�i��iyhhkkkkk]��zOnnnnmmn�qnnZZ~ZZZ~Y�!!r~~Z~Z~~~��cwcsoo~mmmmm~~mn~mm~mmnmm~mm~m~mm~~m~��wwc�m~Z~~ZZq�7!�uZ~ZZZZZnZ�mmnnnn�m��cgkkkkhhyy���ieiiiii����Qa}}}�}}ll�l��}a}lllll�ll��l�ll}}}���������������˭|�v��i��yiyyy��p�[lyi�����������^B^^^x�x�������x������E��qede����������Ž������ī��Ǣ���ū������Ľ������sifdgww�����x������F���x߆�÷���������������������Ѳ���س��������������Τ��������������������������������^A�t��^L�����F��F<����@����FF^^�<FxFF�����@FFx�F����^FF]]Q[f�fiiieeii�iiii�iiyyl�kkgkk���p�nn�nnmml~nZZZ~Z~~Y�!!�~Z~ZQYX~��cwcs~oXommmmmm��n~�~~mmmm~mZ~mZmm~mmZ~\�wcc�m~ZZ~~Yq�!!�q~]~~~ZZZnZ��mmnnnnkY��cnkkgkk�hyiiiye�i�f�ff��P�p}}}����llll}z}}}}l}}�l���ll��qr[b��������ˢˢ�å��v����f�iiii�����fii�����������B�^�F���������x�����t����sedesv��������ı���ı�����ĩ����ı����ı����������dgGv��F�L������^����x��^�^��L��L����޺�������ز�ز�ֳ�јس���������ؼ�������������������������������x��������x��t����@^���<���A��;�;����^�������F���x��x���A���<����]]]p�������i�i�f�eiiiyyh�zkkkg����pOnnnmmml~ZZZ~ZZ~Z~Y�!!Ԑ~~Z~Z~m~��cw�s~mmmmmm~mmmm~m~mmnnmm~~m�~~~~m~~~~\swwc��Z~~~ZY~q�!!�q~~~ZZ~ZZZ~a�~nmnnnOm{�cnggkk��lhyyeiieff�f����a[}U}}}}}l��ll}zl}l}}l�llll���p�p[[[[}�������Ø������������f�������x�������������B��^^<�����������x����E�E����sSdd}w˛������������������Ǳ���������ı��������dedd�Gз�FL����Ԇ����x�Fx����xx�������������������������֘�������������س���������������������������������x�����8:��E?�x�F;�FF�<�A���F����F�F��^<�@������x��xx���^���F�]]]}�����fiiii�f�iiy�hhlpzznnnnY��pOmnnZnmml~ZZZZ~~Z~~�!!v~Z~~]YXm��cwcs]~~~m~mmmm~mmm�mmm~~~~~z~~~~m~~~]��wc���m~ZZZ]~q�7!�Q~~Z~~ZmZ~z�~mmnmnnZѤcnnnn�zpzhhyiyiif�������a}a}}lU}U}}l�l}}}�}}l}}}ll}llh������bi[�ı��������ʵ��R�ѭǒ������FxJ�������`�������^^^����E�t���x���������YdSe�����������ı������������������ı���������ddd_w����A�x����������˷�L�������˷������������������ز��ؘ�ز����������ظ���������������������������������^�B��:8?���@F�A�F�F�^^F��FF�x����;�<��������xx���@@FF��<��]]]}����f�iii���iyyhhSgkz��znnY�аnnmmmmm�qZZZ~~ZZ~qYr!!�~~]q]~~mlscw�s�oY~mmmm~~~mmmmomm~~~~~~~~~~~~~n~Z]�sww�rnOZ~~~]mq�!!�Z~Z~Z~Z~ZZ~z�~mnmnnO~��c�nn���klghlyyyi�����j�all}l�}}z}}}}}}zl}l}}}}l�}�}l�����W�����Ę������JJt����������Ę����բ����f�f�`{���B^Fx���D�����x�A��E������cedel�pi����f����׫���������������ı���������geddVG���xxL����Ԇ���xxx䙵�������ʙ�������������Ѳ����Ѳ�����������������������������������:�����������������߆��;^�x��������xx�F�FxF���F�F������<��^F�F����A��;�xL@��߆^^�]]][���N�y��N��iyylihkllzz��nm�w�O�nmmmm~lZnZ~Z~~~Z~r�!!�Z~~q~]YXlscwcs\o~m~ZmZm~~mmmmmm~~~~~]Y~~Z~~~~~~~]��wccUOn~~]~Qmq�!!�YZ~~Z~ZZZZ~��mmmmmn�~��cn~nnz�zklkkyyyyy����`�[n�l�l�l}}�}}}l}}}}}��}}}l}}}l�[��������ܢ���ī�����J�������L���ȷ���ʒ��f��f�W�{�LL����t����^��F���Ax�E��t�:���r\gdem�����y��������ī��������ױ�������������eddgG����Fx����Ԇ����������������������������������س�����ј����������θι���������������������������������������;�^��@F��x��F��F�F�FF^�����FF�����F���x��x��xx�FF^���FF]]]��i��iHyi��iyhylhkgkkzzznnnm�аmnnmm~mm�~~Z~Z~Z~ZY�!7�]Z~~]]YmzVcw�\\o~om~~m~~mmXm~Y~~Y~ZZY\~Y~~~~~~~Ys]sww�amOZ~qq]]q!!�Yq~Z~Z~~mZqz�m~mmnk~ƹcnnnzzz�kgkhllyhi�����[�}}lllll��lllz}z�}}}}l}}}l}lyU[��������֢层�bb�ibN�||�����L������ű���W��W��{�����L�E�����߆����������8A�ܭ\_dd�Zze�����f����������ı������������y���Ve��kcG���
����������xЙ��LxL�������������ֹ����Ƙ��������Ѳ���������ظ��������������!���������������������^<<<^���FFFF;F���@@���F��F�xAF���<��������A���F�����B�FF]]]pb�iiyyy��iihyhllkkkkzzznnnnmwǗXnmm~mmZl~~~~Z~Z~Z~~q�!!�q~~q~]YmzscwcsoY~Xmo~mmmnmmmYmY~~Y\]~Y~]~~Z~]]]]]K�wcc�mZ~~~]~u!!�YZ~Z~Z~Z~~�znmm~mmnn]ǹc_nnnzzzzkkkkllyhyii���pZ[l}lll�l�llll}��}z}}}}}z}lz��a�������t��ű�����iie�i�b�b��ƫī�����Œ��j������{�L�LLLA�������F��x������:�ߢ��Tddd�Vnf���������������������������y���c���dkVG������BԆ�^�����tE����������������������������������������ϥؼ������������������������������������<��^F���^^����x����F�F���F��������FF�<��;xxx�Ax�xx�x��F<�FF�]]]}����ih�iiiyylyllkgk�zzk�nn_mwЗ~nnmm~mZS��~Z~Z~~q~q�!!�YZ~~Z~~m��cw�s\YX~m~mY~Xmmmmm~~Y~Y\YY]]Y~Y~~]]~]\s�wwcr�~~Z]]Zmr!!�~Z~~Z~Z~�h�zkZmmmmnn]��cgOmnkkzk�kgllhhyyiii�`pa��}�lll�}}lll�l�ll}}l}}}}l}}l}}�������˫ĭ��ffe��eei�ei�����������t�{�|�f�����{�x�xx�F����Ԇ�������������^�����dd�hTm�����������������������f������ccdedd~G����������Ԇ��߷�����E�Dt����������������������������Ѳ������ȹҳ�����������������
������������������F�B<��F��@F������������@���A��^�<^FF����F���A�@����F�<<��F]]Ka��yyyyyi��iyhhhlShhkkk�nmmnmw�mmmmm~m~l��m~Z~Z~YXq�!!�~~Z~Z~o~��cwcs\oYm~o~X~m~mmmmZY]~Y]]Y\Y~~]~]~]]]]��wcc�Z~ZZq~r�!!�Y~~Z~ZZ]�}n~~m~mmn~�vc�mnn�kkklhSllyhly�����}Z�lllllll}l}llz}lll}}}}}}}}ll��l��������ܢ{��fff�����ghhyi����������j�f��f�����j�˷���C���������������������媄�dSeg�������y�f��������������������c�e�kOOww���F�A����Ԇ��F�x��������������D����������������������������٥��ϥޚ��������������

�������������������x���B����F@�@@��A�^�F����x�<����<���������x��x�Axx���F��^<^��]]]a�i�yyy��yyyyh�h�hghgkk��nmmnwˌXnmm~m~~�m��mqZZ~Zqo]�*7�]~ZZ~~mmk��wcs\ommm~Y~mYX~~mYY]]]]]YY]]~]~~]]~]~]ssww�qznZ~ZZZ~�!*!voYq~Z~Zod}�~m~mmmm���nmmn��kkghglllyhyy�y��aa�l�l�lll�l}ll}�ll}l}}z}}l�}l}l���{��t��ŭ�������ii��kghyhhiii��f�ff�f�ff�f���`j��B��C������F����x��������������İc_dHel������������f�f�����������m�c�eeShhcw����^F�B���Ԇ^���xF���t��t��D�t���� ���������������������������ҥ�C�����������������������������������D��F�B��^^�FF�F�^A���xA�;����F
�Ԇ�<^���BFAx�A�A����x��F����F�]]]a�iiiyyiiiiyyhyhlhhhkkk�nmmmmcيXnmmm~mo�a��m~Z~Z~]X]�!!u~ZZ~~nlyc�wcs�~~m~~X~XYY~mm~~]\]]]Y~]YYYY~~]]\]]sswwcs�n~~ZZ��!!!�oY~Z~~Z~��n}m~mmmmOnۅVmmmn��kkhShhhhyyyiyii�}}�l[��ll�}}ll}���l}l}}}}��}}}}l����ũ���ı������i���lghyyyi�iN����f�ffff�����j��{���C�^L�x������x�E��������Ľ��kdd�y�s��i���y�y�����y��������c���eggkwG���ȷ<���������^���xx������D��t��E�  �������Ԙ���������������߆�C�ҹ�������������������������DD�D��F<�<����F���^�x���A������F������<^�^xx�����F��xxxF�F�����]]]ayi�H�yii�Hyyyyye�hgSkk��nm~mcüY_mmmm~~l}~�_~~~]~Qm��!(7�]nY~~mkhccw�s\~nm~Y~Xm~X~~~~YZK\]]]Y~Y�~~~]]]~]]V�wcc\im~~~mYu�(7uo~]~]Z~Zm�Z�nmm~m~nOۅVmmn��kkgghhh�yyyyH�ii��b�l}l}}�lll}zl�}}l�}}a}}l}zz}l��l�������ı�����iii��lhyiiieN�if��f�Wf������W������^��^�x�x�x���x^����E���������Ľr�gd�e�m�cu����������������~ccc���ddg]wG���������޹�����^�����÷��t�����t�  ��������������������������C���Қ������������ޥ�x����E���E����D������^^FF��F��xFF��x���^�x�F�������<���Fx�x�A�x��A�x�xF��B��;^]]]a��eieyyii�eyyyyyhhhhSkk��mmmwÂ~nmmm~m~}}Z~YZZ~~]]~]�!*!�qX~Y~~~~o�wcs�om�o~X~mm~~]~~Y]QK]~]YY]Y�~~~]]]]��ccc\~~~~Y~mY�(!uX~]~~~Z~X~Z[~mmmmmn�զ�nmn��kghShhyyyyy�eii��[�i�l�}�}��ll}}�}}l}l}}}}}}}zzll�����ř�ū������iii���lyi�i��ii������W����W���j��|��^^�x��x��x�����t��������������~cmd�d��~cw�vv�������~�\cccc\���dgg\GG����������������F��������x�^˙�����E�D  �������������������������ҹ��������������������������������D����F�������;���FF���A���F����=:L����Ԇ�����Axx����@AF������^��]]]ai��eie�iiyi�yyyyyhhhhgk��nm_w�ommmmmm~�znmq~~q~~~oY�!!7!��X~]��~~cw�s��Ym~YYmY~m~~~o~]]]]~~]]~]Y]YY]~~]]\�ww�~���]mou�77!ro]~]~Z~qq�n}�mmmmmmmaĦ\mmn�kgglhhyyyyyyiy�����r��}}l}llllll}}�}}}}}}}}}}zz}�y��������竱�������i���li������N��W�f����������j��|�˷^�L����x��������x���������彎w�_d�eeeUswwww���ccwwcc�mdeed�g�cG�����������������x���������x�������E�����E�������������������٘��������������������������������:���D���^<��^�����FF@x�L�^x�A�F�A˚��<FB���������A������F�x��<��^]]Kz����ff���ieie���yyyhhhgk�nm�cȭonmmmmn~�pa��]Z~~]]~Y�!!7(ԐoX~~~Q]�wcs\\]]\~mYmmm~mY\Yq]]~Y]]\�]]KY]Y]]Z]sswwsY]~~mX]�!(!!qX~~]Z~~p��a}qmmmmmmOa�\�n��kShhhyy����e�ei���[��ll�ll��llll}��l�}�}}ll}l}}}����|���tJ۱����f�ii���y���N��W��`����j��������������x�^�xx�Fxt���x��x������x䵙L���׽�c��dgdeefel�ssccc�o_d�ee�ggg��wG����߆����������^F�x�����ʙʙx��䙙����:�����������������������å����������������������������������������F^���^��F��F�@�A�FFF��F^�^��<F^߆��B�x�x����������<��^��]]]U���������iee�iHi�iyhhhgg�nn�cϢ\_mmmmmnz}�׏~~~~Z~~o�!!!(Ԑ�]Y]~]�w�s]\Y]YYY~\YYYoYY]]]]]]��]]]]YY]]~Z]s�ww]qYY]]��!(!7(�Q~~q~~~Z�Ѷ�}mmmmmmmp�wonm�kghhhyyiiyHiei��W��[al}}lll�yllllz}ll�l}}lllzlzzl�����ܵʙ�ū�����{������i����`����������j�����������{�xx��^���������������������xLL@�5��ĭsw�g��d�ef���effffe������\wGw���Ԇ���������������������x�������LxL���Ax��������������������������ؼ��C�����������������x�������������D������<^^F�F�F��FxxA������F���F;�F�^^���^�Fx�A��x�A෷F�A����C��FF�]]]z���j�������iiyhyi�iyyhhgg�nmc��]mmmmmmnzl}�uZ~q~Z~~Y�!!!!!(ԹuQYo��wcsY\\\o�mn\Y\YYo]]]]]~]]ns\]~Z~~]V\~]�sww�oo]�u�7(!!!�Km~~Z~~Z]�|n�nnmmmmmXpm��ghhyy�i�yhyi�ff���jpa�}ll�lll�lll}}}ll}l}l}}}}}}}�b�`�t�t���髒۫�����������������������������������{�LLx��x�t��������Ԇ�������LL^�x����zcwcqdddgg��������dd���cwGc�����^^B�������Ԇ�^��F����^���������A�F��^�^�������������������������ӆ�������������������������������^���^^�F��FF����x��xF���F�xF�F�F�^��B^��F�xx�A���F^�Fx����^��]]]a�������`��Ni�i�hiie���dyl��_c���mmmmmmnlla�uOZ~~qqZY�!!!!7(CӅ��cwcs]YYoYY]YY]]~]Y]\~]]~Z~Z~~~~~~~~\]]�K��w\��u��%(!!!!!�]Y~q~~~ZK��Zy�mmmmmmX��wX�klhyd�i�eiylyii������pul}�l�lllyllll}��l}}ll}}zaqp}���`�����J���ǭ{��ѫְ�����jj����������������������������xL����������x���������^^��x��ֽ�׮cGwc\nzkz���dgO��cwGGcN����߆��C�B���ԥ^xxF��������Lxxx������xxFF�F<����˥���������������������������������������������������������B<�^�AF������Ax�F���<���^^^^^��^���FFF�x����F�x���������]]]a���`�������iyiyhiiieie�y[p�_c�Ш_mmmmmm�yr�rZ~omZZZYu77!!!7!�-�ucw�s]oYYY~oK]K\KYY]~]]ZqYY~~~~~mm~]~]Y]�sww�v��-,-77!!!7C�P~Z~~Yn\���ynmmmmm_X��wm��[[�eieeiiyli�i�`����pal}lll�l�l�ll}�l}lll}ll}[zp}}[�[�{�ūŒ��{��{�{|�ː����������������{��������������J���L����������Էx��������x�xF��߷����������scwGGwwwwwwGGGGGw��������߆�������C�^�xx���������x�xL������F��;�^�<����ҥ����������<��ѳ����������������������������������D���߆������FF�@�xx�����A������F���^<B�����F�FxAF<��E�C������]]]z�j��W��j��W��iyyi���eee����y�̫�_mmmmom�yU��Xmq��s�]u!!(7(63�(3!!�cw�s\Z~\o�oY]YY]Y]YY~�]]K]~~m~mm~~]YYYY]swwu�*,+7!(!7ځus���~O�֌l�~m~mmm_o��why���eie����yii�f�W�����a�}llllllll}���}}l}}llll}l}}}}r�u���b�{���N������й�`������������������������������t���L�L�������������x�����F��^^�^^÷��������Ķΰu������u����۳����������Ȇ���ԆԆ^x��������������൙�A�F�@���;�A������������߆�������ކ����������Ȇ�����������������E�����DD�����^^F�FFFF��A���F�Ax��^F�;����߆;�@��F���^�^���A�����<���]]Qp������������f��f�f�i�}��p����vՁ_mm~mm~�z��Y����usu(!7060.%!!!��w��~Z]\]o~~\\\\]Y�]Y]]K]K~ZZY~~~~~]KY~�sww���1�0!(7(!�������Yq��n�~Xmmm~mX��su�r��}}���fff���W������al}ll�ll�ll����}lll}}lll}l}}}}a�����r�p[���N�`�j�ʗ�������������������������������JD��x������^x���������������^�^�����^߷�����������������������^�x�������������<�F����������L����EL�x���x@��<C�<^@F�����������Æ�ј��������������������x�����������������������^^FF��FFxx���x����@��F���F���xF�FFF��F�^;@���A���F�<]]Yp������������������}��qqZq��wwv�~Xmmmmmm��Z����'()!τ�!!!�6�cw�s�]�]�oo~YYYKYYKY]\]q]K]qZ~~~Y�]\]~Y\sww��!1-.!76*!*v���(+'�u�p�~mm~mmmo��ww��qZqqq�z��������������a}}llllllll��}�llll}z}l}l}zz}}}Upau�s�s�qU�����������j����jj�����j����������������JDDE�x���������������E�E������^^^B����^��<5���������������������������������F�x����x�����t�뵙�����<���^^;��������������������������������������������������������������D������^FFFFF����Ax����F�����^@F�F��<�@�������F^��������CӚ�F��]]]Ub�������j�������ї}�aaz�Y}�w��~mm~Xm~m~z~\��*))/̎��13M7��wcsKs\YoX~Xoo]YIK\K]�]~]]��]qZ~YZ]]YY~]swwu6-3%61,!����.+)(s�Y�ommXmm_o��ww�z]y�a����������������al}�ll}�llllll}ll}}}}lll}}zp�}}}[}PKKsss�s�up�����Ê�j����������������������������JDDE䷷������䙙��tt�������������������÷���������߆����Æ�������������F�F����x�����x�˙��t���xF^^<��<<^�������������������������������������x����������������������������߆�^^F���;��A�����^^��F��^^�^��F��F7<���^<�����Ԛ�^F��]]]Z����������������b���}}��Y~�wwϫ~XmmmmXX~��m��(+)-�us�-�0%6/!!C�w�s]\]]~~Y�K\\K\\K\]\]Y~~]]]Z~Z~Y~~ZnZ]sww�6�%,�s�-+)+)�~o�zmmXmXmXo�Єwv�Y��}}��b�ʳ���������}l}l}}l�ll��l�lllla}}z}}}z}l��}}}aq]QQQK��s��u����À�j�`�����j��������������������J���L����L�������D����^�^���F����å������Ȇ��������ݷ������<��6�����������Ȇ<��x��������������L����A�^^<F��A;^���;��������������������������������������������������������D�����䆆����FF;�F��F�������;;�����FB��@FF��F�;FFF�^�;����CӚ���^�]]YZ������������{��``��i�}�Z��w��pmmmXXmmmml�~~�+'(.څ��-�,,7070��wcs\\�YoYY\\\\]\K]\YYY~~Zn]\YZZZ~Zn~~~]scwv60!-7�s��.+'(�~�zXXmXmmmX~��ww�aZ���N��||����������b[�l�ll��ll}}lll�l[l}ll}}z}}}}}}}zZ]]]]]QQQQQ���uu����j�����`�������W������������j�JD���xxxL����������������������xx�x��BBB�Bå�����������Æ߆�^��C��������������Fx��E��������������^�xx^^����x<<�A@�^���;���������������������������<����x��������������������������^F��@FF�@��F�����F�F�;F�5�^�FF���Fxx�F��^��C�Ӻ��<�]]Z}i������������t�||��``������wβo_mm~�mXm~��oYZ�1)(⅁C**66!,-�7�cwcsss\]]]]]\\K]]�Y~oo~mXYn~]~~YZmm~Zm~�sww�!!!-!!7rs�())�]ZX��z�mm�~~mOm�ǅw��}����|{���ŵ�������b}�ll}lal}l}}}lllll}}lll}za}��}}}}Z]Y]]]]YQQPPPUp��v����������f�����W���j��������j��� �