SYS9000/04--,,,,"-"""$"-,4449997900,,,,4l�܂-.��zy��#8v��im�G!:���Hf�K���G 7+���I fUs��S�oF=���-���~Y==I=H\mmldSSHSQSYWWWYSEMHHEEEEECEESQGYhl_��~YhhlSSEECGGG?<<<<<===<74<<=IIQSSSEE@9999E~�ޟ-&��zW�lv��izoF+���So�K���G +:+���IGWi��Sy{F)=���4���~h==EES\pllSldSSHWWWLWYMEMHEEEEEEEEESQIQqq_r�qlYllqllhYYoaWLWWQQSYYSIIIQYYhllllldSSSSSS~�ަ)��zo��#i��nzW3~��Su�U���G 4F	+���I UUP��H t�F97=���4���~hIGGISlmmllllSSSSYYWWYSEEHEEEEEEEEEQIIWhq_��phhqlq~llqqqoaWYWYYhYlYSQYIQhYl~lldldldSSSy�ޘ +��z~�|#*v��iEG3���SW�K !���C 3<-���QG<g��E o�o=���/W��~lIIIIS\llldylSShYYWYYYSEEEEEEEEEEI=CIIWhq_p�{qhqq{l{qqq{aaWYYYhYhYlYSSSYSSlllShqhqldSS~�ކ%��n���##|��n4G+���M	FWF %���= 4<+���IQ<i��E o�W=���-	�Ɏ~YQIIEShlldllldSlhSYWYYSEEEEEEECEEEC=IQSY\_p�qoaoqq{�@2m�ooYolh\b\llSShSSSSlldS�22m�SdS~��:!+�ڀ���2z��n3U-~��MKF?!%���= 3:-���IzE"8i��; o�F=���/���~YIQIIQSlbll~lSdllYShYSQEEEEQIE=EIQC=ILYYYYp�qxoqqqq�;,n�qqoqhlhVhllhVSbSSSllSS�H2m�SSd~��4+��z"���;2���i4f:~��HF:3+���= -F$���I�S61l��; o}F=���,6���~YIIIEESS\lwyllllldSYYSEEE9EYYE9EQH=EIQYQYQh��uoo�qq�¢��qqqqlllbllldhdYdSddddS����ySdl~��G!%��zo��SB���ml�<{��M:G+:���= -F+���Q�l0o��;h�:;���/0���~SIIICESSSlqwlddldSShYSIEEEQYWI=EQIEEGIYQQQYq�xooqqw����plqqq{llllllllldYdYldldl���SSll���z!%��z"���,;���i��W/${��P?U+���9 3U0���Soo)
Y��6 ~�<I���@4���~YIIIECSQYlwpwlSdlSSlSSSEEESYYECIQSIIEIQQQQWhq�uoqq~���pm\qqlqlllqlqlllSdYdlllllSldSddl~��y %��zu��0H���ml�{y/q��POK+���9 ?U-���SWu)~��6h�b	H���4@���~YIQIIEQSSqlwldSdSShhSSSEEEYYYIEEQYSSCESQQQYqxuooqqlmyml\\qlq{llllhllllSSdSdllllSdlSSll~��)��z"o��!���mW�~y/���P�{3+���9 GF7»�SUW ���6 o�GS���C@���~YIIQIIIQhlqllbSSSSS\SSSCEISYYIEQShSSEEQHQIY��xoaqqShldSYYlll~lllllllllldldlllyylllddll~�ޘ��z��f���mU�~y/���X��3���9 d?E˻�SUU���8W}4	V���P7���~hIQIIQSQYhllb\SSSSSbSSQEEEQYYIQSSllQESEQQQo{�ooYq�~~��~�~��������������������������������y4��z#��W���mUe<  ���`QW<!~��9 YU?���VUU���BWo:V���S<���~lIWIIQIYllllSbSQSSSYSQI=EEQYYQISYllSSMSSSWhq�oaY�����������������������������������������S:��z"��o,���n?W-���gE�E,-y��E {� G���VWFW��Dou:V�ƮS4����lQYQIYShqlqlSSQEQSQSSSQ=CIISYQQYhlldSSSSSSYq�qY{�����������������������������������������/3��z���0#���m4U3	+���i��M'"���H~�$	C���VW<V��P��hg�Ȭd4�Ο�lSYIQYSYlllhSIEISQIhYSIEIIQSYQQYllllldSSSYhq{qh��������ª��������ڼ�������˰���������	3��z���R8h��m4U$+���i��g**���H��+y���d�l0	P��g���Eg�ͮO4�ǟ�{YYYYhhYh{lSQIQEISYYYSSISYSYYYYhlwmllllSlll{qhl��ί�����׊�����ڬ����z�ھz�����V�$F��z���@/g��y:W!+���s���68���MW�4/���gV�6P��g#���,Vg�ȮE-����~YoohqqhlqqbSEIIQSShYShYYqlhYhqhqlwllllbhqoq{Yh���G���݋;���z����g��ڝ����P��qB����ґP�43��z�}�Y��m	FU$	3���v�˸cB���S?ob-���gzy#&v��i#���i�i�ͺM/����{q�;;m�ql{llQQIQHWh\hY�55g�YYoql{llllldh�V@g�Yh���4����i2z��R|���8��׍v���|1���Nc����z6~W$+��z"y�qq��y	FU"=���v�˼�����S:WzF���g|�N.v��i#�˾|�i�ϻVV�Ο�~q�02m�qqqqhSIQLYYlh\h�M;m�hYhqhqlylldhV�S;m�YY~��5����Ds��.v���v1`��cj���c���Pi|�ؿX2WG %��zI�Yd��m	GW-i���|&�˺�sͻ�SW��Wh���g��sT���i#�ɬ��s�ϿP@�Ο�~q�¢��ql~llQYQYYhhhY\�¢�~YYoqhllllllSh�¢��SS{��1v���D|��.c���c1N��iX���T|��>8v�ٿR*�l ��z"QWm'6���m	W<7*s���v&�ˮTd���V����g���X��ic���i�ˬzI|�ؿN9�����p�����{qqqlYQWYooYhll����lhYholllyllSlh����{YSq��H����Dc��>v��c.j��;T���c���c8v�ٿR*�� 	��zYl�>>���mU-5#N��؉&�ƺc�ƻ�V���Vg���g��Pc���i��|BH|�ϿN6����������~�{{qlYYYooohoqp���z~lhYqlqlylllSll~��{YY~��i|���>>��.T��c&v��V`���c&���cDv�ٻR*��9�ڀQ��NN���m	U4"*R��̉&���|����V�Ɲ5����R��0"���i��g2c|�ؿR2�ɟ���������������������������������������������������Rv���D1��#Nv��T*v��zz���c*�Ƭi>�ѿR�~d@�ՀQy�M0���p	UU *i��و&��������V��P2H���g��$,���i�o�gv�ؿRB�����������������������������µ�����������������������8���D>v�2Hv��T*T��zz���c*���D6|�ϾR��P0��z<�����m	oo!	,���|&�˻z����d��)8d���X��P/���i~qS"Pv�ؿiP������������������������������������������������������P����Dc��1�k��T.v�˝���gz��`6�پN*��B,�Հ:�h	���p}}3	+��؉*�ɼS����V��6N����Xz�;y���i��QPsv�ؿv`����������������������������ڢ��˟����Ο��ޯ������g����Dv��8ji��T2|�Ƌ���Z6��|H��ؿR*�mB4�ՀGoU���l}�U 3��ى&��U3U���V���Nw���PlS2����i���ccv�Ͽ|`����ި���ˊ�˼�¾����ڿ����z���{����q�������쑀�΁Rn���Dc��8vT��T&���gP|��g8��RE|�ٿN*�E �ՀUoG	���m}�U!:��؉&��+%o���V{�y/F���RzVHR���i���vcv�ػ|g�����I��ݮP��qV����g��Ŭ����B���z���ڀC��o9l���VE��z>R���Dc��6cT��R2���PRv��g@��;P|�ؿR�7�ՀetWW��mf�U%l���|��-F���VWK	g���R�7*P���