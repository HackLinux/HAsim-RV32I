�ǳU��&�JDjD��"�Պ�92�J'o���E��Xq�sya������b&�Նe�Y|��u�,G��+�EJ�uy���tc)n+�F?7!y�r��u�@^�B� ��C���XX�B蘱z�����[�wQ��E��^���o�Еa�cU@��1l'�T5�����N�(���`uwG�.=~��e��3���>���~�Mz���A�^�o���JG�H�Ͱ{�PЧCkK�i5��3�B�>� "m\��
Eٙ��������U���5���u���qgh���Y_3� �YAxo1��e�A���ʔ���O��F
���?�����nzLUxy�8��>����[��ŷ���?c�Ή�w���p�V������E����c`�U�+���~{��t��F���R�h�Uٚⵆ0�8Al��S��]/��l���D݆^�]	0��g�e+���=߅^��'y2���WB�У�-���ԁ�i�6��8�����*��	3��ג�������K��g�G�c���G�ْ�l��o������ܦ݇#q���.f���UxD�.^�)9BJf~��t|����\�j����>\5��6���ܦ����^���gΓ�*`?�����4�/lg��-��[Xv�Aa{�:��KR�?�c7i��l_�00޻�Em�l66A�G�p򧔿ɦ�%MՅ�dc#���ü��R���ݣ.w����-�m>�:D��9�7u���ӢL=�ѩ�-R=����$t#7pF�LM����QBt��*}�lx�/B�Y �ދ��ߒT;2����f	�ŵ�I����ԎNd�7wɺm�0�@�P��v�ѳ��ӧ����[��lua.	���=}�{Lo����6:�éS�穐[��P��<��3���/�"H�_��U~�䔧d���O4bh����B�lr,v�u��/.��&��h9��� _�J��'�p�|����ԊQ�հ���h#c�`^a��r��i��rp0j���� pl�s��h����Թo�Z�Yl�ҩ���8 ���t����J�eh�=�s�����qv�ʅ�{R/� �E�W�̔��T��w���Xt���j�J��H�p�̹�4�\���	����9汿z��ܢS�R�ΕJ�W8�ٔJ���r���S�	�G���Dͧ�(���w`�`V�&�K�n��6�"���cȕ㝙ظq"�.��Ν⺦ �%O}gK[2�򬬸�n^�a�ǻ��i1�4�<'ü��2گT�Δ��6��JH���^BX���Y��!}�/�蒕�Ũ(�ZL�]|���^*wZv]CᄙƇVQ�'%��c��3�g�lUAΔg�BZ4<-!�
kZ���%�����Y����n�?���x�'6J�QwMɢW�Ъ�%CU��9Sv�*��ӡJ�O�~M��v<��\gT-N𦛚3�VϦ�*x�[�z�P�(x��*�}tH<l��UR�'���/����Z<���oFEr�t���@cb�}g��7(U�S�ElMɮ���x�V4��u;���}BZ=/���xA�PÜ�΍�gQ����v(7F��PἝ���I. p|�X=�l�qT�A�����$���.S�|]�g
7 �^Cɗ.�n���#=������c���ud��i����r���>z#���g����)Dիg��q��/��$�d`��H��rl���MK��(�w�Q<6|G�a�����a�@B�ɤ���GR(��OH�$�	|k~Him�P]����X`tJ�V�Oh�� �Sҏ���Yj|L�Qw�\}6����W.�0�x��Qm����my�mw<x�3s�wQ��}�;�|x�z�s��e3����LoD�=���*�h217����e|TP��#���0,��Ȱ��D��;47r�jX�ݹ��Ga��Ҫ����#��[�0��@~!���(GwU-��L�$����|�w�ؼ���ʛ��(HbI�~��?�c^�%�� &�Q��_X$)��s�q��O��/|�e!��e�;������Z�E�$��.�����0�E_	����e����|���.��,��&����ʯ�{��l���P�5�����~�����ؔa~,�i� h\�NY��V��
���q切� ���uM��x�����)J|G�^�|�]��z��н�~J����j��1��A�*�)��ʞ��o���P���\\�"�0�Ek*ˣ@L�ĝ�tD�w�*� ?�Y��)&UL	�Hh�#�o�1\BM<Ml���?<��Ek��O �?����@�9IDG^A�+�",)7/�A+l=�'d��KT,D����s\����h���t���/B4����Kp�u��|�O�aT����C��7Q�z\�����=��&��EW�d%Ī��+C}�]p!y{Cף[n�ׂL;���N�g�`�z!��o7(�'^zG=_~���c����*��s�t� �����;'w|���vs�%��(ծ^&n�U&�_�ǹ�$����:fh2a#��b��}T���vd�t�B>���� 	F8'�D㟑�RR��'Cc��As��v%g���xc��' ��f����D=�<��¼j��-�7�Ծ��<ѿ�Qj��/,���t1:�
����U�[�*�&�d�˥�_����S�j��lrN~܅ /�M���c/��s�OW#	|�kt�$Q��N��6O.6_#��X�G����Pz�m��'K�!y��[���ЃU��{�"]�R�ڌ��@�(�q�SXj-r�@yz��HA�O�x2��p���	*ZJނ�'Eǖ	iاqu����	;���ם0!��S���;|'��E(O-I�e�`�}��Z�	�nC|=@��
���� m�r�<*@~&/7��σod\�x��ѽ��E6"}�5}K �A	�)�xKYɠo+H7�/�~�`�T#D�Y�����H���%�L!�$jh"\>i	z�ݺF�J�h8�06q�ܤ�탇3��d���G�r�QT��[���vR�f��6ʈUN԰U��^���ժ����;�>�g��Պ/l�T�U6ݐ!O:	���Y�����'������+�%!K�A�����r�r�O��i1�F���/w�I|�k�b�v�N��I�����Dɉ^Q�3<DL��oDD��H��y衋�㏢��A�eL�
~����?'~z,ǹ����y������ݼ�_�n�\zԇ/kι���p���g��!++��}&��V`+������UD ���'~��;w;^%���8�s�5�%L��R�-4*�d"��-B�q�����H��>�E�rαd�UmXRO�dE�Y?KZT�~��-�[�Bg)'x*R���P���ĥ�a�,P|�Kп!�`�U�$0��@��0�£��0���)�Wq�����,�����J:Ert� x������%[�bܷ���V�@���݊��E\B�CȟF�����'w��vr��o�>��{�����ݾ'�K��9�m�;�'�\V��s� �_̋�+�⮝��*T���As���}ֻ�|����.���3�l��pxq/��|.~��/����0(B#�_�[��� ��h�
��T@��H.���#��1�ͯ���i	��6|����iv��#u����FZxf1E�q��)SNݺ_=�EQo��)�$hm�~�M��E��{#ʫy��c:�(p��H�h �XGj����,�}p�=|9��5]�{<5�j�"�[���qP;�|�����Wl{�PD"��h&��� �-GRi@��������v�K�%y`g�?h���㩭����b�`a�{���˃��?��C��7�}�j�ǐ�c8��d���QR�.����.:��ټ�w��b�_^�䛽��`�=o}�o1�:]t�b- �*\7�~@��u����k�����Tr/{��R�e�O�&S�^���7$���&�tZ�������H��u��˸؇�:�b2;Ѵcj�&�p��b��y�X��1ݐf���ERz�V�z4�3�|K�A+��i`��d�H�k�k�d���p��HsS�4�u�a��ux�����������π@?�`���[�n&�{M�XrCP��ᚳ�[���\��������o�r�LA���m����e�$�C}�����3��>����0�>�#�����28�*�b5�V���w*/�H�P���X̛����r��7�դ3��'�k&�q&�NW�Q���?��(�8��~b	ܙd�vO���&Ljͧ]�w������Y�9'w,I�36���D!�H�hM��G�g7kQu�-�c���nA?c��2w
 �3\C)������e=��3̢�=��\̴��8�s���$6Y	)��4�[��T�f�g1V'g��b�A[�ps0���l�U��]��o�Rwj�3�8"�\=&�����I4j�zH��^NӁD_웲v�&���[|�c�8dR��zTw�"ʘUl��$f�����3?��I�X����{֔i#�;; K�#����3P"&՚����A��r䮂p��)ǋҁu���Y��� �O����0Hl�_%�Iv���	eU�R|���y��x=�P��*O�4➫��uꒀe-nN��5���:��q�����5ul�M�c-�T=��TR�T��f��m���&A�J�ˉ8"������� G��z���#���o�]4?Bf�2;��:4!�'���)k�k���`����_L����f1���p�>�T\ٷn��׃*��\H���`)��DS�[t��.��]�}�����:�SB@V{��_��郉/b�>��_"��+��N�ݛJ(-��g�����4Jơ	��Ň���QOB��:\�J:�ܝX|�!4�ڠ$h#���kNݮ޿˭O0��=�t��^Z�S�������R���Y���!�q(��R��h{���_=}uk�73�Vj�A4�%��b��r'��]f����M�xG�a[Ivm�o�K�*F,��:�=�Xa�+5�x�<�f�u=_�}��*H7]m]����^ZRd�l�F�W4I���������-��˳�)(�kF��OЌ�џ�[�o�a~|���/,�4<̩�%gZ�n��t����A���J�B�v��
�8�s9�ʹ�G��+%d�}Ȩ��w�*_�b]o�&JI��q�.��Uѯ{ ���k��;��2�j���(e��|���V2���D�XzS��e82໖j���Mr�oqၮ�,�fAWsiV�y 0�����r�x��NW�e��n�f�X��җ�K�jh��*/����\R�HZy��Y�\��*�3�+gmŋP�YG��oQ�_}�Cͷ5t'�7_r�͢�w���BQikh��-�#<��D�Y4�f���2��U�>'W.�]P?ä��5���f��KbD�i�V�.����󜁡�`h9���aj�}A�ةi${P��Îz�LY��V|�k��p�}��<���2Q�8r7�~������ӵ{^�7�����G< �vs�����p%��Gqqy@��8�׎�^�L`/�,e�/����lO�|�+�۽Ǣ��t���}�1���>��q��p���L��+bdh�!��E�s���x�l'I���F��X���(To�ȉCz�F���qY���1TyZ���c-�+M#mH��2��/eZt~���4�6w�W� ̣�����w)�G8U�����M]ӝ�CZ��_b���HEΗ��2��
(!��xS�\���W;��i�O�F���@�e~<�f�4��l�dq��U�p�$/=?%6ݖ�j%�	G����Х����+qWBؔl�!!.g8G����W�^�?#�OBA}����Z��%��)�ȿ�X�z���b�wR/.9��������o�M���fT�Ix;gi�+����y"��K�o���$�hܶg��[0�̫�8�E�Eu��Y��e�!�(�[�S{a;�AP���j{=���g0���3�/HO�:��0�ܻ!9j�
��嵆�	^���0�׀�<\p�"��o{��[��g���0��Ԯ��Έ���*��ןw�ٿWN�*��p�>�zm쉈
 ��ǖ�}zElx�x���nF>��Ȕ��,>^s����Y�ʐ	\�3�a���@ҧ�}�<-�-�>�Ua����.�[
b��٤�9%�\�^��^���=N)f���{��{�XP(�/�v�2��@�Z��	�Z���X��?�����>���_�������vE�7����"2t�����m�cj�<�6:eL]ѐ�~1hO§��3{t��:��(E���.��~ya!��u��G�x�Jy(��꼳�eR���|g��$����f�74�M���G@��6�_�s{\E6���N��.t�)�u��;{��߲��h/��-i/��)iB�6%�/N
j�**��uMt��K��v��q��e/^\dN��?�S���Ն@�O����ou�5oߒ�K�t8�hA�n�G���a���f�nCrq����)F�Yh��Ղ�T�X��S�ǈ`�Y�p^�[L}p�eK��%O5x6s5������V��PP�Ȧ>{0�e�0l��:]�~��߹a��Pq��w��ktl���`�K˸�A�F�=K�+���=@n^<�@�$�������
��<�St�D=��n�R:cld4�@�7�M֓\��a�`�P�����?a(jh(b(�=;�jY;h����狊G�#�JC%Ǯ��9��T� ��.f[\B.T��;�I!���W'��w6�s(�q��|ړH#~�HE�Q����~��q��1����b�aP�$XT,=$���r\|eق�ۯ��?�`�ַ֠G�����y��wɯ�]{lѫB��_
솦� ��;���+(��"��&b
_&r5]@��W7c�Ѝ��������L����c@"�j�;?K�@��̥����+�˄oE��J=����i�o�Tl�{=��"b�^�����i�fw����Y*PԵ�z�x�D���Z��F�s�9��|h._h��敁RF�p�nNB�O��{���˸���[0�zО}�$����އC3k?����|��/e>$|��<�khN�L1�w�1��}n��,��=�>+&�U�[�\�GA(O��� 3�KQ݂��krƫ��k�Q	���k�}����߆�}�kV��;�(O�q�o	��`�?�;3H�ļ�3u���x�	�?A��  �[@M������l�Q8��!yH�sO}g1C���!���QR'	��Ωv#>�_?�n��s'^��O�	c���A��o{�KWO)Or���Am�~�/�"e�o������"@w �I=��j5c��72�ŕ��/9��Qp�ȇ�N`pzUPw>|���]��.7�m�϶�lW��v��%��$<>i��,�{�M%������>���xt��h�uY���N��L�&�t�f�Oa�n�c�JU���-zb��J�a��ze*�'�8 F���.3�yl�st���cKo�MƮ���"��F�◿�}����X�Iخ9{^����ko৔ې=|���糟��`eRa<��\���]����~x�¹�igh��'�i	��;?�C��>���S�BD:v�cߵ���,������ܝ����� �jJwpH�yP�>���I�;�h�/a�00�����(�^)��@���y~��.]��n��g��#�ݎ}�'ʢW��$){f�m�BQ��9�[����ݕa=���w`\��噻�w�Y�<��59�&2��h�q2�/��F��Ɉ��4����Ҋ�?>�cGK2F3H�$��T!�E�!K���Co���O��؁��6Ce�h���)Bgƿ8�3�ɔ����G?����!�����7YC.�t� _��2�1x���J��'���}�NL
���xD�"ڶb������)��������B	��b{�f�I���T���D��@^{����٣�%�\գ,L����D��$'��p�����q&g�����N�ߙE��۽|5|%"��۹|����E�ftidݻ�%O�!��!�0{� HP�AI:�R#%7�oC�P�|e��KSr���|�3�D�����z%K�k{���G�� �(6Y�q�J�����粞q�0���`K�n�`]�^i�o/KQ�d���	nmB�w���.��h�k�F�R�7��8�xꞟ����\;�ݨG���8n�ɯ�Eo��o�w���;��/�����n��o���=�S�/��C�_� ӪXv�H��߷zX��*����d��Bm�N�6��&.i�B��B�����)��u�=���P4�"��X��S����x`�wʔ�?�t�u�}�-{Zƿ,�>+�۟ߓ��KO�T�o�*[U�s�����TǜƟ�ص%�� ���x�b<���&xs��ޕ6�o��yZ!�+'��_I�9��������JZ���?��	em��00҆6չ5,�i�m�&;���=�6�|F�-'���C���S6���"<�n�o6+*�05(��~�)I^���˥��Dou��Ӏw�7�R���u
M�/I����fK�O	]��	���`0'*\:Mp��&�&��T����n�ʠ�R�Lmخe� ���q%'�^��`,�����	��Lq_3`g��sj��0��i/g:�B��L��J��������jp2-Ы����_7����Q��Pu���%�H��[ApE*F�'W������*�U��~���hָ��c�vA�,����"	.؍Q̶�{z(��<���h?z>�sn�H5$~�]=��]��=�j=~��_b-?��?B���maz����ݕ|��vy������\��(��a��ˀ�F�q.���]�!:{A�;F,�+��	�+�;A*�n_���d�������{��v>��u��B ���Z�㡐o�qo��C�x�=,�T3��W�����Pz& 
 ]���`&4��*��U�9I��	���ED�OJ�[��?8]xOHSp$Qmw&��B�%�q�M��	�������?��,4A%G�f��/��[�dK���	{���)S�b����ܳ��>o�a9A��(Aܛ������"�ܽ����{�{g�0�X�
?R#������n+I�o�����I"�Kl���� wu]� HU��=�=�g������7�s?�T� ��-׺Y�ut��� ?�#�����4ph��Rc@��~V�����2��	j8~�>���H��廽�:.8q�{n������MX�V��o��h�)���q�Q��?�n��3�#��-�x��V�d\��K����=]�%P̘�ӠJ���J�J�JO�<�x�w"t|���]Bo��4�每��©xR$��:��D�)��pLod�U�l��~_��8���I%�3�S�H�k���VMrgA�
��ҍ� Bp�N����4 �b�+���B�;WӻN��~[�B�؉7:8b�6>�n�Ż=��>3=`qu��һ�h�.�`%������I���A��a�~-qW��[~��gkj���\d���M]�I{�U�Jo�b"�f� ���9D��J�$z���!U E˽��$ 3����Vk���-�J�)��˺����͐��\�y��v��r�	�8�SA���Y���y%G�u˦n�� ��굥0[�_��#X��1b�gb�O'8(옻y/����?^p��8ÀE>%�}U2�;_WÖ��IOO��f~��|��X'a_(H84���n��Z�D~Qs:}��W�D��0[�&�og����JN�`�����"`/���L��Xc�W%�F���.I���;���B/s㇂�G��ԾE���4cf���q��G������X׏?
(΅���_#�;y����8I5���y��Fd&P�����\%��U��,^��L��U���$�����M��|�>�3�(0a?]Q�k��e�~��Q��\Q�0����9u���	*WN-ChF��i���{��/Wf��!s�|��i�}E�bt����m-��o��z:������V��|�K����3F��m���{{;����7�Η��P�ە���<peu�Ό+}�A��w�zN�.�����p�_y��߃o=�+��; �	f�~�ҡ���*��(�C�}d�s���cŢ���,�9ʖ+��.2ބ���h�%���iƵ��2C_@�u+<A��j�=R�_�C��C��gj��ŗ%J��5 R�����0~v9djx*&~��}�|NO�3�>e�v�`cu�Q�Rz���ϧ����)<�� �U@sfa�{�f��(��d�Ԥ�)��~������Gu�ď17a��׷'���Kb������}��β�̥U�ޙ�1�M�}���r�N�M����9�=��&�1��:ĸ��l����q�*wT�|'����v8:�t�N] Ӷn�G/[����8�R�`���8u�R�5�%�" �~�s��g��x�8��?Lnq(7Y�O _o�6�]���}8�|!�p��V�Ħ�� ���Wa�-BX�G*+:�����*�`�8�~M�b�����;�����uE�0�R\�]���!�@E��O���c~6�=A_����F:�&v�2X������%�z�/ܽ���$T]K@KՇ�ڜ��B��@'d�h��}�?$��'{�þp���#�}�A4�[���{N��Q*@DR\g[���z��׊j�K�{�5B�����v��^��d۸ۼ��(��:�A�u@+s��D��gC����`S��)��X����4S
��'s�ȃ+v^D��K��v��;Lk�R���{�n�T�?��-��^1��z�~@��Y1�"$8{��2�D(���PU�0�
�WS�nr�g�Q�G$;#�F�e �Ik��Y���0��hl���7�9M>�7�MKH=��A���&�_>Uw�?�;�b�I�ΏW�2����K)|ya!x�{�/�9���^Kބ�E�r�~�~r
[:l�5r�&����!0@ltqe\��eN��wV�l{]�IP3/�_�Et�~}~>�͵��7���N�h�cұ���m"�I���_���b���}@��5�ܧ���`x��� +����$�vu
�M31ҭhMS0�����0�N�Tg.<��3ü���t��c�di�ƅ�s|إWX*Հl�Z��T��%�%�'���;=�,��럃�t�S'n~`@�b�'c�EQ�;M1h�� ]���e W�HO�o�l�HO�Dc��!I��2��`�NZ�f\ڎW�D�sQ6_��qӥs���n�k_���g��q�>x�s�g�e�gq��c��2�s�_P��9���R�^_ԛ�[���f�s[Z g���Z�ng>��d�dh�u�{_ �v�]`Y�8�W���B����]��i���SXS�ɨ�P���
�Y퇽��:X.���=I�&�nX��_����3Wd�9�c��G�x�����
�"�k�����58���zk��j�]�IF *ܪ��D�k�ДИУ�S��6$���N�;ԕU���%�`��'a����Ą�k[��mDL��(/�y���5�s��_OܱtAoH6 M0��zۋB���T|k>�qi�R)����BY�n��h)Κjz�G�������LK��#nC�H�l�Ĭ���ޱ׍�~�T �앓R�*�7Q��x�ĸU���XqU!�ӁNRTm�(��ݪ��8�
m�|eU6~Y��B�����'\s�m�޼P���P7����+ʩ�Μ_:��M��2	)�}*J��^����(b0Χ��w6�n�ۖa� �w���-6��]��nc�RA%�`�O��Z��gZ?��8q��v����Pu�����L�W-�W�=⣯�<�Տ�8�&!x��PV�VQ��p|kv�60�T��b���|��rw�ߐ�r��OM�j�|c�_md��;s�jN��vCI|NiI&�YPۅ��cj@j���m���$������p	���^���t$�a�&x�S�uk�����B�����̛�b���?�/�O#G^�߮��0NǮ8��%��=GV�����H��n4�CL�~<�(�?�Y��h�x<$1�"�B�/
6fTɞ���ybңϲxw�[����@H�_'�PTaam!;�>��D�#$ecO�ݑ��������&�ꃗ=R�p@wDsjj��S^��e���4G��.�F��8��/����7�n[
�W�7' F��{]ɂ��p���Q��;��k���k�o��}X�a����Ḁܑ�J�� �ܓ4��$����5v����X�g�� �D/����40T�2q��x��?�\&H)�6ך{���y��H�)+�A�>�#���l+V��Ƣ;~��pk <�ǭh�(�C�R��l
����D?�D�:!�����r�GlsAL{)���-�h?Y���4목	�)��pL(��6<R��Bڢ�b�]B��b�0f #�k��~���[>��4�I���!K��(!`~��M3e�N���?:��~�|�<+��u��/b#� a�{j�e���](�Ρ�H5�㈄�BCm�^'��I�vй�����Z��>��dp���i�B�"�id�+J �=ѬE!aa�V(�ZX͓i"�,h�-�+�-~�B��-�?)��VN�قzρ����u�ruf��ƨ�u��l��uy�/��`s���i7�Ҝx�a�v��~��E�e?e,��;�c�
��T����%N��Gx<U��l�X��>�A����%b�8��>B 4ɂt��cc	{Y?x�9Ϣ�Ay]��7d6)C�.#(G�G��R�&�����W�
��}�:���gU,��� >�!��y���Ao\����X�������]�|~OYO<�FK� Ci���#�k��|���݄�>{��]�]�+1����t�44 �w�L`b��"��6��|��L����-_��u�6O�t� ����۩b3`��GqK#��(
pI	��.9L��mЬ��g����R���S��`�R��X���+ �^���ӗ���po�7g�G���j�C��*�7�w������y8	hW�e�-�}�B������+6��q�(�� ��4c����Ͻ���<j�|�/>|��`��nL4�.�X`���NG��$�w
2�f	��������y��o���3���	>cZ*aɌ�Z���R�>X�
6�|=��fpu%�����Co��k�s�q���}?"����c͒%2F���o�_ ��G���x��!���i�dx�FSV������(���.��Sx�����v�5E>is��g�E<�p��"��8��]tb,�9 k-s��+�P�ɬ7r�!w�C�