�"+�g�����������-=��6lK�^�ؽ�a�&ؿ�	���?�C��\]�[��OMצ�SäN&�߲�Wٓ7�MIn��Ъ�iS�	�ԣֆ���:�>�Xe��^<�9Hx�k�������S�d��'"��fԯ�)4n�z{Si�}�AS� hm)]V�"qǆ5�$���B���ѺS�{��h8*W=��uc� ��>�Yп����0��ۚt�9��Eƞ�k�r;i��@�"/)U[��O�P:�إLQEN���,β�i4i<Zx�n� �A�"��#��b����e����;�M�96��q,̊W��,4� �M�0Z�ڇI����;�n5OC�>Bxj���D��n�1��#��ORd���k�����#�d&X��M��:2�]� _7H�f����EٌܫH����NIhMq8gV�괇TVq�޴��� �Ӱ�V�����h!� �; ����Ή�z����i�!1p����(�K(�<��r��Ru8le��P����ȳ��Oϐ�_3b���g�;\?)�c
����ƴ�M�D�6;�@��,�1��K�� !�O�(�#NV���&��02��gO��c�?�=���G���8�"&��T�aL�{Zq�ڹ�����Q�L^)������ȑ�y2�8Ӯ����ٍ+`?���< �o3x6�}�ap萅Θ�62��Z7%. }�h��S3�R��s �����Q\��5��E6���cX���x���WU�#����I�Wd߉�q˘P�P���e28ſ�I���_C�eT�66�/��o�z3�ϠƜj�4�`�;@9c��+FT0���k��\�{�σϫD��[q�4cZGc�<��Pv��^<�ǹ�%A��4v���,��l)mk֝�2�hY�FX�<����k<��DH鮃@����uPtơ/�1Q�(N�P��kS'�jw�7?¾���ڧ7��tEU���}͑��z.��'ED"<涓NDՏ�ʮ�M҇h�qA�Ϙ�ڨ�OlZ�:>h�x�C\+vA"�d^h� �=/e���52Lf�k��gC������������k��ʴ�^�,z�qFE4Lx�0�������L3��P_�翇CE�Sғ߾�f�u��ݚ�s繏�#d�P�H�\�2��td�D�O�&��9�U�T�<WH�"�4!�+�~R�J�6�h��W,M������ل�X.��r�Ѣ�Z���/L�|E��ǲ�_ҏ�� Q����mD]��um��^��!���q��o�;i����}�!,	B0M��Ds������k����=�N������ѯᏔ���q����jlĸ�D����F��j�N��J��WQG�R��M�V�9/;���a_�·ޯ8�|��Y�l�d�T�x�b�`����^�C�f9n�N���a
#7k�gj�|~�������rL˝��Q��*nJ}�x�YX���[��65�&A\��6;�(��c~'��''�?�ys ��~�.?��-uTìSj�M'2<Ff��G�8|�k�[k|P���A;}F8�F^�Զ۠5�����G��V{���I;+�Cqx��9����v��Ϟ�s��8�j繶x��x��l��4�ތ�����f ֯�-&�8� T�ފǹ��o`�à���14�H�Ů��^RȘ�ݽ|[.j�tЏ|�I&��+,��fF�����y�>���3�Xi���I�DG���se a���v/P���>�7��0�,JS�dIm:x�r���u:���A�����j��q�� X�ʼ�T}����Q��pi�S��ܡ�����v��HҰª��*i���B[J}�щP��.�e����{/�4��IN_���u)����NE$�*���ezS�X�Fmʹw;	z/��Ư'�Ew����'������+�֠�3��*P]�,'�Ud�{92��͊�g�>8�y�'H�Q0t��SڡS���V�P�@;9dߍ��kO�K7�
�r'�@g�Z=|��;��� ѾS��������p2�2,tZ��O.�'
.�h3m:�$����7��Qk0i=;~���]:,�y�k
�8��v����ԍ)����n��8�Y�T���K��lP(x�[�������!�����N�$8��Cc��R\��p�V饗ӿ�������>����o����A��p�J��߿���
Ĳ��'��Gm,3+���:/�wơ�n\���n�jW��t����!���Ѹ&�;c�B��$U�[՗��v�S����'�S�x'D�6��hiԙ0���s{[n@U��:���V3�٦�=�G �c�)*��le@|���NKv�f����$�BO	����<-�K �§�Bw%\#j�ʗ����m5DW�����؋)Zw���A-��c	�g��V�B�ʌ�J�N�)/WյO���tH)N���q�X���N��xI�b�:5���Ņ!��#uv���^����R�~Xp�rU~d$�C0�w
��.p׏
A$K����*���uoKA�0>�/����c.���(����	���A��\�ܝ�(����@{)�F�`�D>۵���r�tL�d��xȥ����;��W|:���s�6ш��lq*5)%��.حK���:Ug��1b����bSa����ӱ�ܣ:�ӱ�X���p��2���%3�J�{��aߴ�<�����z�x#�R������2��|2���C��VRJ,Ҫ��IM����s@��z �Mˍ�
u
=]F�w�T��?�k'ԫO�������U�A�l�W:\R5͕W��y��1ݸuKw�N\� a�����IN����?-�T��[|-tL	��B&9��V$��+��bEm����]EU'�����D[�{)�z�JZkV!�!�R��T�L:��UP���P̅��=���i��X!�N`��E��`��m�C0�0�xj�R�K�iO�9G�%�4箔 �ԗ@�3�зI�`�	�>�x�I�)�M4�/���:����@������*�/*ߩ��ݞPt�J�n������u�Ns�� 2;�T��^R�� ����u�uD2���~t>�4�x�n�!Z���n.���� w����x+���n��S�vk�W@n�2s6]��p�]z�$
͆���#�Zw�����z�4x=1�-6�*�ր0,&�%WC�`�ܺ������싵%��ۺt��z̓��c+7{�$s��n������)���y����=WZ�h�j��d�.���+؜u������Tp����ṟ��j�`�yH����o�7��<�H>�z�����A�P�Z~ �팮�R�����l�J��P\"�x|������)4=c����&��˪�ЎV��g�-�uƦ5�I �ĳ�ٙ���1���#�������[;�l\�����*3�_z'���#Ta�r��k���5I8wwsD>��Z�5o>Q2:�ƀH~*ý�����o�K�/[@Yඎ�[���*2t�R�=�k�n��!��Jy&I4��"2�y��<��k��id�,<*xk�`�s+|vCV���o*B5��OI���kF%G�5�u�쯞���p�H!����j���(u�$�y`�Z~
m��ϴS7�����y��ゲQ��fZ��7�S�zBL�С�OW\x̖��CcFG3���Wa�w��2\<"�O��ަ�3��8�*���s�>K��x�1�َD6f�W]��h"��/4h�7]�@����4/o`��4�o`���c_��qo4�t�;�`����3(.+Ýn<� L�(��xTG?Y�Oj	������i��eh��J!!0��7�m-mBlD*u���f��>��0"�NfL����!�[�/M��b}lDa)�j�"���CVz��ܛ7�"]�e��'7���7E��,��$箌���w�5z����kY�X�6�yY��O ��c���,����yJJ0��۫�%�&�����Q���6�	�`�Z%�5�:�������������=��tsl<-%�O����3����x5ۖБGȑ��@���������w��'�4�h�y���qN:.Ev�;j}'-�Za"q�E���`�W�u�~5p�f� �iW��9��hB�@8l�-R�?�S�=<�_l,��� ^��N/ݼ��	i�����']qgݦ��L�_�2SA�����6�93���R����o��Y�dn���)�3T��Qg5�Oϸ�KB�3;�r XQ�牢eRWr�� V��gHaï�3l���<N��}���#�x
�ַk*v\���et}�O�w{"=x��|�{�$cJË�K"B�o�P3F�p�jW�@sש�Xq�Ap����Wb�� y#���ލ�³�mi�����q͜���Ė��5����a~�FD侖�..����-t���Шq���#���R���d�:Ռy��{�հQ�{4*��g$E#ޖT"�_Uz�R����rc4��]d<�{aT���=�O�[OP����ը�)ɠ�ð���K2�,���kr"�V��z����A����x�Ÿ���mɴC){x�*�F���x�DE��\n=��r��eG�
}�e����0*+�emԎqU�wٹ�3�#�1��c�D%�fuS {ƥ������N���g[����Wt]39��������	E��slA�j<�� ��"~3C���i����B���b]�]c}����t�a�Z��b�Mqc�1H�����++�xMlE��dU[��[�7�mv���@~.-AfH�[\���^������~���X#��]�$�!k�Jp%�����]�:�{��ѵ�[+��5E���5��w��ʸ/�@�*C�@E��|3p.%���3���Wo]q*�,L$~< ��S��oI;�:��䔒s(a�wb��b��[Wt��X���:*oy@��Ld���=�îFn)�K�%��B���'��#�-6�jQ�˫�[�9y������ڍ2=́�q�6+wR��
�	�za��%��ч+���P� o��JeW%�&����xf��5f�l)�S���%:�Cc�BQW�$����K��ͮ0����������}�y���