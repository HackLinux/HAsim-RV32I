���Q�B�@�M�U���E�M�d�    ��]� ���������U��j�h��' d�    Pd�%    Q��|SVW�e���t����E��M�U�Uߋ�t����M߈��t����$  �E�    �UR��t�����M  ���t��������j j �p�
 �E�������t����M�d�    _^[��]� ��������U���<�MċEċH�M�U��E�M�M��U+U����B��tG�MċQ�U�E�E��M+M����A�х�t&�M��M  �EċH�M؋U؋�EԋM�Uԉ�E�K�E+E���@�����A�х�t&�E�EЍM�����MЉM�U�R�E�P�M���F  ���M�U��E��]� ������U����M��M��/O  �M��A�U��B�@Q�M��Q�E��H�J�U��B�E��M��U��B��M��Q�E��H�J�U��B    ��]����������������U��j�h��' d�    Pd�%    ��   ��X����E�����}� v�E���T����
ǅT���   ��T�������X���;JwUj �M��� h�, ��H
 ��Ph�, �M���s���E�    �E�P�M��>O���E��E�X/( �E� hT�- �M�Q�Y�
 j �UR��X����HQ�UR��X����HQ��X����O  �E���X����B����X����A��X����E;Bu4��X����Q�E��B��X����Q�U��E��M����X����B�M��H�e�U��t4�E�M����X����B�E��M��U;u��X����H�M��U��E���)�M�U��Q��X����H�U;Qu��X����H�U��Q�E��E�M�Q�BP���m  �M�Q�B�E��M�U��A;��   �M�Q�B�H�M�U�BP��u,�M�Q�BP�E�@P�M�Q�B�@P �M�Q�B�E��R�M�Q�E�;Bu�M�Q�U�E�P��X����8K  �M�Q�BP�E�H�Q�BP �E�H�QR��X����K  �   �E�H�Q��t�����t�����M�U�BP��u,�M�Q�BP�E�@P�M�Q�B�@P �M�Q�B�E��]�M�Q��p�����p����M�;u�U�B�E�M�Q��X����5K  �U�B�@P�M�Q�B�@P �M�Q�BP��X����YJ  ������X����Q�B�@P�M�U���E�M�d�    ��]� ���������U����M�E�H�Q�U��E�H�M��U��BQ��u8�MQ�M�����0��3҅�����t�M��Q�U���E��E��M���U�뽋E���]� ������U��j�h��' d�    Pd�%    Q��  ��?3 3E�E�SVW�e���`����EP�M���q���E�    �M��Q�M���q���E��E�   ��`����z uǅ\���    � ��`�����`����@+A��8   ����\�����\����U��} u�u  ǅT���$I���T��� v��T�����X����
ǅX���   ��`����y uǅT���    �"��`�����`����J+H����8   ����T�����X���+�T���;Us��`����p�����  ��`����x uǅP���    � ��`�����`����A+B��8   ����P�����P���U9U��  ǅ���$I������ v�������L����
ǅL���   �M��鋕L���+�;U�sǅH���    ��E���M�ȉ�H�����H����U���`����x uǅD���    � ��`�����`����A+B��8   ����D�����D���U9U�sD��`����x uǅ@���    � ��`�����`����A+B��8   ����@�����@���U�U��E�k�8P��I	 ���E��M��M��E��U�RQ�ĉe������������U�Q�ĉe��� �����`����Q������� �����������`����h  ��<�����<����U��E�������������������������R��`���P�M�Q�UR������P�Dw  ���Mk�8�U�щU��E�PQ�̉e���������`����B�������������������Q�ĉe��������������U���`�����g  �   �E��������M����������������������������������������������������8������������;�����t%�������?���3Ƀ���t������R�F>
 ��뾋E�P�8>
 ��j j �8�
 �E�   ��`����y uǅ8���    �"��`�����`����J+H����8   ����8����U�8����U��`����x ��   ��`����Q��������`����H���������������������������������������������������������������������������8������������;�����t%�������/���3�����t������Q�6=
 ��뾋�`�����`����J+H����8   ����������`����B������������Q��<
 ���U�k�8�E��`����A�Uk�8�E��`����A��`����E��B�  ��`����Q�������������E��E�+E��8   ��;E�"  �Uk�8�E�PQ�̉e���������`����B�������������������Q�ĉe��������������U���`����Ve  �E���`����H��p�����p����U��E�+E��8   ���U+Љ�d�����`����H��`�����`�����h�����n�����o�����o���Q��`���R�E�P��d���Q��h���R��s  ���   �Ek�8��`���A��H����Uk�8�E�D�����H�����P�����D�����L�����^�����_���