�W���'�Kj��0���£9��w�A@9������0e��naI��$�`kY�;���/ܴ�Z�����k�ȳ0��V�X�3�s_�_��8ٶRx:p_���𮭠�̬�l-K� k�� 9Y�9w4�^]�?�cT�s�I���v���h�wRtt=af�X�0����p	44b��V)��<0�q^�@�֌��˙P�{��\b1@dA�)Z�>00��8�4(��@�q�G�d�����sl����	�wp�	ӽ�-&>�eY(�9NA�CJN���h��b-�ۀ/)Dԁ��=9H�SW
�������)�I֞}A�]��g��S��!~
��	N�������o��l�VbZ8 ,K�+IK; �����ǁ1���:GD�����3]�*s��Ɔ��86W�I���}F  �D_�.P狏A$g��C4��0eL�J�'EE`J���#�Bk��c8���!�H�����S�QgE
� ���I
���R��T����"ݤso�����5�=	vK��<؅8�8�B*<��G���� ��7@�na\H=Z��wn�E�P*����s��0�����T/|�1����k��! �eM�T��y�_��os�N�"��/�VW���m�� ci��l�~�u�-`|�56�+<)��E��]3rS1J��+�h�5�;�kg=���~)��o�ل] [|��#��N�?� ��#oS��M��]�@�qh&��ڴ�}�����v�=O���9���x�a��V��?���~i��;V �i�fݷ�>���M-D{5�9vce(C9�B��CԚ��+�e�.�&���A�SlBnHq���S
��M��\Yy "�F��s""�Ը���C�9��hFi�<��Q�3T���;��ߦC�L��� ��ox`�������Ҁ;K�IC��
���'V\3��vP[\���d��A�j�_��g�E~D�`s/d�+K�s�_l�sٲӀl�� ����:�O����T���1r�(��������a��T ��,
�� 
��r_Y:��Ƅ�����[� <@9�"��H��{�R�y���K�Ez�e�$`A�$�M'�R-t�6[g8 K,>��4��⢅��7���I�9x�yN~^(���W�B�^J���/�"��5�k�:;��3h�k���%�}A�vu�J���C�W�\��KY���������Q7����Q�(�[��$N��F��7�.��vB�`�2$���B�!����� �J̕������nI���ݹT�2�f�o��b�2#&yw������q�y� uh`A�'��R0z����h)����Pv�Y]�0�yǪOY���E���is_x�|_���_��Z���~�N ��:�!;[H�6س
V��w�o������f����ף����kL���m���?��%@�{PiH�U�M�X����0W��F����Q�Q�,�~�v���ޙ��X˲1 ���TmL���C��n�+ �7|���dy�y�;J�j��J��)��JE���g�t2�����<�ʝ�b��Vo#�,L�������'�l��#�µ�K����
(Sb��F�iC�||`�$K1�թK��CD~��:5S��_��x�7��( ������<Qo��)�S���7_Z��,ړ�"��x�TJ���N$�6t62�ϩ������I��췗�h�_߽�6�mc);?���z^,��Z�vr���R��䨷Aլ|�L���*�:�����{Z������~�����h�\��5"��m^�ɯ��b�G�ltr�FfB9&p3���&`kX	�4:�&(��%�&��oi�LAɢ�Pc� iF.O�ɶcqz��4d�Uib��$���}��S��>��W�Z�\�����ӣ�W<ѤkC�'=6<jAv?k��$C,���Y;1ɲ�X�zH�ǵ��G�?���UB�[���Q\]�M{D�R�X6B�i.o}Vh[Y���A\1RvW���Q��T$D]�����Z𛄪�),�Џ����C�Ɩ�RJ�!�6ס?��KXi��?��S��:ؽ�i�<�펀�^�n%�BJ�	�]�6m�e&��.H�ҵ�4�[iw�-屸����I�H[����e��>�Y�tW�-��2�k(TL�����;B�� �S���h�M�<R�/��PO��}r���t+���5]�y����y*�`y���n���|����Ƿ���2�,�Ω�r�%(��o��Y,�J1���-��C�Xt��� ���v�>��$̈����Z_���,J��.Y�ן0o*�㸑�%�d����R�=�F,Μ���otU�܏i6����/E�����폿x\�*:W�Ⳋڭ������'HBX�F�i�Vf����1z�J����p!Eq�|�/�0m���۴V����e�V,0�����2V�`646��c�"/$�r��6Sk$�%��n_��SDD*��������Y�NV��BꚄ���y�X^
�Gjc��J��:�+��m�p������]�.l����]���6}���~���*��|��U�۵E�ҋU�$f�A;��f�\�n*3f=�Wۚǿ�絎8���9����u���>�Iw:~���Y�$�?]ſ�Q����B����R F���`"�