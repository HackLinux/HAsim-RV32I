��|���1�\kAe�@/�y������ڹq$�Q��es婖���Ps���I���i�Y������˸���]��Bēl��1��Ԓ�u���}�`����T�6�����0����֬.GL4���i���M[ּ9Z�I� �GGq|Z��r�`�Zcr�g��(����0���VA&��6��ͨ^G�.�PsE��(�o���p�X����a�ÒG�E|���ƀ��0D17�E?7,���g�#0N�����c����-J\�#JP��oTA"i�̗�Ug �e�n
|`��^W�d�YΨ�(�6c�o���(��V�J���"��'�]�o@UxH����f��x͐� �ma*cG�*;0�s�h�y^ח�0���)@xD�'��rB�A�'`x��u$դ�wr��(�i%v���i�bk����B+1�7�@E�r�Or���м�IF%7�nA�ba�eu�n���]�.�l�@���%9�G����7��5�dG�yթ/���r�f�	��NJ_�/J\Ѳ���$0�!F�'�td��m�C��~0���D57�0��[��Lz����>��,�1@md���A����s"k9͑��Hb�u�2w�(�t����!˖�̐�v��/������RШ��U֮���ݕh�tD��wX���d�se.q�y|��y�ɡl���>uÐ��(�9��d0��0��%��57�Gdߖtc���$3��ԶuC�vt��q����b�c�A�T_��B31R�SF��yu���7|�����!�\W*i�n�$�Q��o+gg��2����4����3��.f��[��X�Si�tD� ˗����ﹹ���YVeMT֥�����I�����`�\V=p��'׻���|�?0���A���ud�^��ES�QgE(6�~󯠼�׻�>�B��!�nGDֶuc&��t�U��B01jE�ܟd�w�|���|��f=l���nH-�Z��&%7�Fz��b{���鶚C90a�FG��t�w���G{�z�#�R�6�@�}�w},��8����C0�o@5g{�̯B�yk(̑�)C	0gD���g0�i�.��������F �޳V���C0E��vP��n�u�!I���T�R�5B
1ʡ�����~��ˮq��}*p���׻��Xy�0F��ͯ��琌\D!7��o,A���Z֧1�FAj �n���3�AJc�۶�+���X֡B0�*�"�j����[�|����-���~�T��C60��PG,#
G463Cs9���I��䚘L�ce�^a�^����\���=u�������2�zA�©��t���@'1b~Ҩ����hY�_ѽ�xU6�?@m~x` }�������C�[�ệ�����#ejq����6�[х�7��@�7�Y@��Gr�Q��F�(%s��pY��C)0ը&GTC�̀sŤ~��h~
_�}Q�FC?1�CF��j*G,wAu�� �hruȆ��T%������0r�����(��X�Y�����D��E�>����B$0�B 0�I
D(6�����g���&���Z5�m��7��-�Ey��P��nt�7%���z�6�ґtĆ����jl��^�'���*��Է�j,���#���jlT<�M�;1(���}��%	�"7tbj��/7p����[��T�7��k�m ���tF�D6���t��o��Q�^��Ֆ6���Ic�������0s�Ѱnza3|��ȩ�(��'��S�Z�4.潐_|e�i��%Ϩ|�?��GUס�'[GD!��S��1��u�u�9м�ҧY�WФ�&\Fz5F���Wr*��S�0���T㐰���e!]����w\�a�[ѫ�y ��\G<6���g<Պ�j7��&���~��%s{2�%��x�����a2�L��i�t���xj*�J��w�M�df�[Z��[�\���S
Uѵ�%s�{˯�"��e9ɱ�F`���Z ���&f�j�?�t����m���G�b���A~d������z�Y����oP���/0��or�7.1��F$7�;�Vj�4�[@] �% ��;�3.dF#�s��ʩ��1f$Bt��G�i�>��|%70�7F�a���sїr�(6�~>���KY��E6�{7�`���<-�G��Duۯ�Ks���$�.ɩ��XP�x� ��TЖ�Xйx?0�x/0�x��x��0�̫t�Q3�<A"�Isq�� �nD�hՑ}�Ů�d+}����
^� �nGs��YW��x�8F@F�FEtd�g��qP��C1z�QF3z.�A�t����o�m%i+���1���A$0��m{@h
@1 ����1�	G<6��Ԃ�bL۵�_�e�W���YЉѱ��超�t��Q�$���' hTQ�����1��^Cl%�����
ZѢ��cY�z �u�׻1׺!7�=7�-�����ؑA}AR��Ft�ׅ_�������7��v��Щ����,6{�"A
�>A
�.A��6Ar{c�P��P�%!1+-6!�6�6G��j���n������0,����A
�$1���ğs"����iW�-1��E(6;�nA�zï`����Fq߯`��y7�x����ӡ#/0�įŀr��þR�F��t��%t���̨�Y�(��\�քCpT��Cv�!��os�y�x0�����owrE����1�F6�}���@s%��G�(ۂ0���D-7l�m@��/͂���ފ]Ѳ�2�FC���/s�I'}�y�Bś����+f���*30�}��)��.���������Ӯ�g�)��"�h����ud�_�T�7�^Q��������G7�E(7�:��������r��#�l��;4��y�.c(̑�DS�GH�:s�o���R4�=0�B0U�.G���ڸ����*�͏�Z�T�Y5��cs��y.�����Zփ�F 6#xï�z������/q� 7�D7����ž��g�Ʃ�n������j��=@O�1����2�F�� �
���1�1�����,c��п���W����������Ʈ٦����t���֔�~�FW3�
�o���]��/s>�0�
A*"֬u� ��r��P�x��W1��ׂ��t���9KT�	���EtQ�J�ۅ%=6�yj��aW�z5�\G$�^u�-k�_���>
^яYV6����6�@=�@}q@x��wUї�AYA����/�.�~x�V����d��a�o&��t��������t��yt�p� �n3�.�"�ϖt�g{�/�.t�I����ݧ!0�$E���"�C��/���K����ࠠIqf��eF%z.��n�Bd��P1ͅ������4�e{���|���O��q��I�Ȱ�e�сu�n��a���-�,㑌��@ZW�'5���<�x3�����̯�%�ʩ�cĜ��oE7�[������J!n��5��D��Xr�j��>tC��r��J��Ϩb��hs��ч��u��������h��=���ż�Ѵ���j2����4�x��A_��1���1� 1���!@e�����Z4ԁ�����瑨��%���v��"iC1���@%��ݾ�<�]�:�뤩�A����Ȇ��6B&1���mt�p��A"�j��:���G�\��7��C06�C�M��&�
�#6���h��K�T�5�A�n�{֣���v��fa;�Wп1��C�.�3#A�o��{
���
����x�3NfB���g�E��
'`��bCa�8B@{����iT8�1 �:gE�%�r� �/�������pFJTѴE07dx����͓�U��]�XʭjA�ɡ7���e��6/b�螋��2ֽ~K^�GE6�z��`����x�[���d���K�F�i��0���u@����uĕ��/�~��K�_ַ6�k��{خ��
�	1j���/y�'e�(p�x1������uğ��o���1��ӯ~Ab����t�4׸�N�1�YFCz��'�wr�v��5�X�z�i8C��w�C1r�z��)��W�B>0��!���uø���q�WЧ�����QЮ�ѷ��:p����@�:�:���@6@��u@ä��u�P�x٦�1��åזu����h���J^ш���|��L����~
i	� B��_s�!���kftd�8���̭1@���r�r��@���=�*0�$��prE�fuj'~�o�D�@�XrE�������"����s"�x�i=ֽ�2Kn�bШ�"c�pY։2 +7��ցt����/�[hft�q1����0���%@E��(P���y�\��F0F��rB�7s�-�͐�nC1ּic���u��U�#�3
SѪ0���E!7̯y@��د�����t#+s����>LR�|hau��@�Y�#�o���e׃���3.=6A4�,G���v_�9��7��i-o2�i�c�vF������_�l����	��e�`��;�W湧~�z����(`�����֭����i.v�~�4D�r� c}[�p����}�!G����A
��pZ��n���gKRЃD��b�!ձu��{���dvA:,����
�/:7�cowr�f1̊���ר��a1��G �6���Gdږt�7�߹ַ���D��Gr��a��-թ\G����Xr%�_�n!��yQ���Q�A%%20%y2Gd���v�n�csg�i��h��ַ��Rƫ�`#���/�]�Rf�BtPE17L�Y@aE77�i�&����s���'����eu����M�X׸�j��&���'��z
�!�yu�=P���4����k��`��s��ƯЦ���ɵN�Fo?���vM����1��<�$�drB�?r�c���>6��t6���� ���@�6zrG��l@�(�������]��E7�����lf��h�����V� 6��H6��ܙ�G'7�D37�_@��#r��.̗�C�2� A�{��@�f`�n7��'T��6��SZ����G7&0����v� ��Ǯt�7������`d�i����UA-A���Ȇ)�HZБ�c��ݹu�ש��͋%6g�(�/�ͯ����DFr����(�i�U�=��O�m��=�E��n�tG�)�.ʩq)�	1&�4�@%�+E�t$���/�N�o4��xF=���c�[�G�
���{�n����P��xʨ!�%�$7�E'7��¯`��n1�y3���q!�7,�@%"�q^�1�l����se�&�Z֍B00g$7�D'7�2�v��c3|��o5�7Ћn�sE��s��b�)�h�F`w�f�X֎�