��~��~�}~�~~~}}�~|������~|~��}}�������~��}~~|������~{�}}~��||~�����}�~}�}�|����}}�������~|�}��}��}|z}������~��|~��z}��}~���������}{��}��}y���{��}��}}��}�����|x�}~~��}~��~|��||}~���|��}~�z}��~|���}�{�~���~��}|���}z}��}z���~}���~�}���}���|��|~}~��zv���~}����{{��|z�~~�����}����}���~z�~��z~��}�}��x|�~~��~������~|}���|}�����|��|}�}~���}}��}�����{��~}���}{z��~y|��}~���z|}���}x{��{|����~�|}��}��}y��|}����~{~��|}}�}��}��}}���z����z���}~����z����~~��}{~���~}���{{��~���{~��~}{����}~���~~~���}�~�}|�~��|~��|��~�����~}�|����~�}��|��~��}����}~��|�~~��}���������}~~�~}~���z��|~~���}|��|}���}~~~����~��~�|}����|����~|��z��|����~��||��~~���~~��~~����~�}~����~���~��}���}|����{|��~�����~��~��{{��~}��~���~��}|��}����}�����~~�~~~~~�}~����}~��~~���}�}�}���~}���|����~�~�{��}���|�|��|~�~��}}��~��~�~�}~~��~�~~��}}~�|~����}���������|~}��}��}~��}��~~��}z�|}�~���~~��}���}}~�~~~��~���~���{|��{~���~��~~|~��~}��~~��}��������~�~}�}~}��~��~���~~��~}�}~������}��~~~�������������~~�~~�~�����������~��~�~|�|}��~~��~~��}}����~�~��}��}~��~��������~��~�������������~~���~����������������~�����������������������������������������~��������������������������������~�����~�~��~������������������������������������������������������������������������������������������������������������������������������������������������������~~~}}}|||{{|{zzz{zz{{{|||~������������������������~zuplida^\[ZZ\^_dhkouz}��������������������������zihcb\SSUXWSYcfdgqwvwz~}{�}}�~y{|x|��z�����������������|rinkRMXWOJL[^SXdimiiuvxxs|�|y���u��������������������{rY]hSBDNUG=Rd\V^mxqkv~�}x~��~y~��u����������̵��������tn^\X?EF?B>INRR_dfnou{}������~���������è��ӿ������}nZMPE;<;=@DNRV`jmmsw~�{��������}�������ͱ���ð����{vhaG;F:532ADDO\ejou}|��������}�{wx�������չ���ʴ���|tu^D36C5()4EHP]hqs����������}xslnr������������ĵ���mlaK9&/2'03<KNav~���������|}utojib`i�����������̹���xbSD4)$*+&/=M^gy����������xpg`_^`c_`e�����������͵�s_VN>-,;@LZcs��������|ztcXRNQU]hllvz����������Ʋ�xYM>;FID<16J\w����������ycPLPRVXQNPWk�����������ϫ����yaSA06ER\_aijo��������qfccZUQHCDKYeoz����������ӻ�����vfZF6<L\iqz�|y��������n\NIKQXVOLMQ[m�����������ٻ�|tnlpleVC@JYm�������������rXB68GYelie_\gx���������Ƿ���qe_Z\VOVajr�����������tdZMB>CQ^djrqqs{�������Ͳ�wnnpoicXKFPf}�������������lVGBDO`pzyslfgm}�����ʹ���{{xumcXQS]p�������|xz����vi]VX_eimnkheipy������Ŵ��sollihga^ap�������|qhedmz����{utvrh^Z\`eoy�������ǵ�}eZWX]fmqsw��������scXTW`mz����������mXKIMWdq{}{x}�����Ū�]HDM_t������������x`OJP^t������}������re][ap����|tnlmv�������~qqx����|tllt������{pknw~����~wv{�������~yxvvrqrstuy�������~tt|�������vqsx}����}yy������}tnnsy�����||}���zutw|������xkc_am~������}|�����wqnq|�����uoov����}xvy�����~wqpu~������{x{���|wux~������{wwz~����||~������|yx}����yqnnu������xpms~�����xtv}�����xpnr{�����|vsu|�����{xx~�����}wtv{�����zxy}����{zz}�����~zyz}�����~|{|~����}|}�����~|||~�����~||}����~}|}~�����~}}~�����~~�����~}~�����~~~����~~~����~~������~~������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������pddhs�����uhbl�����xmlw����ohmy�����tlnt�����uaW`r�����qhmt~���whm������bKFXt�����ta\iy���~zz�����{rmo|����zkejr{���ypprtvxy���¼�vC4;Z���ɧ�pWN^rz}�������sc[i����nTENe|���hXXes������ɲ�t@(8^���ڲ}hfEE]kgs������ePi����{ZRgsxx�|dbppn��nbfp����ڢ? #�����>39G{����zyz��|^\_`myi_bnw���zqtps�����ӳ�N09^���ÝqXUe~���taXXds||rkjmoqpkmsy����������ӽ�a?=c���ào_ejv��ujjppptmTObkq���qimrt�������ȱ�s]Yl������}nhiklnu}}undYLSit{�qfak|��������í�u^ct������pd\QWl����u\GANfz���mcagt��������ŧ~kddx��¹��`HGTl����r\K>F`{���xfSRcv���������{nbez������ZJGSl����o[LEOk}��}ocZYl������û�|jck���Ŭ�jHFYk����n`VMI]y���xg[Zbm����������pdhx��ʮ�rKCUj���p\UID`���qb]`fm~����ƿ��ket��Ʊ�|\KXg~���r`WRFUq����w_Y^gz��������xibg��ϴ��]EOev���zi`H9Pp~���o^XWXo�����}dY_���Ī�_HLaw���i\N>Kk����ucY`dn��������oa_s�Ƽ��aGJa|���}i\H=Sn}���w`Yabj����ʽ�ue^d��°�y\JXt����vfUCE\x���}lcglmz���ʿ��ca_|�����`WTez���|k[DJ_o{~yotrhm����Ǭ�e`e�����s_[bv||�|ofUIXcku{��xssii����׿�q`Vk�����fPObz~��}jUGO]ev�~|yurgq���̻�vcd����~fZ[jx�{smYHPZbr}��yvujg����̯�jdn�����r_\ds}yvsnhTJX`i{�zupvusz����Ĭ�mku�����q_ao{~woie[UX^`hqt}{xujn����ukm�����ucahw�{mlne\X^ZYkwx||xukn���������������}yssuqhnpmiZX[Xartvzwyuqu���������������wxzzzrcfjjmcdc]bortsryxw�~��������������usz��vkcahkjkjgdhqtvwxvt{�����������������|}}{uqkkmqoljjoquzyxyxx}��������������������~}zxxwuvwxxyz{|~|yy|���}~������������������~~}~~~�������������������������������������������~~}}~~~~~}}~~~~~~�������������������~~}}}}}~~~~~~~~~����������������������~~~~~~~~~~~����������������������~~~~~~~~~~~~���������������������~~~~~~~~~~~~~~���������������������~~~~~~~~���������������������������������������������������������������������������������������������}mh}��}tv���}y|���yw|���zy~���|}�������|~}���z{z���|}~�}�����|us{�������}tsv~����yws}v{v{}}wx{�~�������vx���{{y���}uz��~xv�~�{�|�����|x�x�w�~�~y{��|�w����}x�x��w�u�o�y{�j�u��y|y���xzx�z�k��z�m�v�|�w�u�t�x�~�}~|���|�x�}�w�}~�w�r�}�~�����|�z�y�y���|���z���y�y�~}���z�w�x�z�y�x��}}�z�y�z�~�z�{�z�|��~�{�|��}�y�z�{�z�~�}}�~��}�|�|�~���|�{�}�|��~��}�|�}�|�}�z�y��}�}��~�|�|�}��~���{~�~�}�~�}���}�|�~�}�}�}�}�}�|�~��}�{�}�{�|�~�~��~�}~�~�~�~�}�}�~�������~�{�|�}�~��~�|�}�~�~��~�}����~��}�}���~����|�~�~�~�}�}�y�{�}}�~�{������~�~~���{�}�~�|�}�~�}�|�~���z�{�z�z�y�|�}�|�~�y�}��|�~��z�z�~�}���|�{��{�|���}�x�z��w�y��}~~��y�}��}�|�}�{��|~z��x�x�~~�~�}�x����x�{��{~�}�x�{}}}{w~~}���{���|�z����y�x�w�x���~}~��}~z��|z��|�r��|���r�r�s~��w���}}~��{�z�}�~}�|��~�v��r�o�o}xxpy{k{n~wrn�w�~���������������������wqohmacbcd_fcghfnlqnvs|ny������������������xv_`Z^_`Ybivtyz{��zsokpie\`]_b_^����������¿����ptf\JEKJRZXcs~������uslf^\TPYVZZd����������ľ���wbbVE;:LLS\^t��������yvrlaPTFQTRSY_��������ٹ�Ĺ�~pg[X<5:RKN[bv��������|z|maOTOOVHP[mf�Íſ���ݱ�����oePW=8ILPKant���������zyu^SSSKLPNYcrj�ɍ�����ঽ���wp\YOA6ITJWXkz����������}ygWVTJMKOR\jgr�ʤ�����˼�©�zvhZZD:EPPJZ_k������������tdbZSNKIQXZehty�ғ�۾��Ŷ����x�oZ`HAMQNFYaax~~����������lpm[UUSOZa]dpx~{�Ä�Ϯ�ĺ�������tfoVIYYOJ[VZoqp}���������y~yjqlp`rx]}vd�{}�~����������������yiikcWZ\O_h]hrq{{�������|�v�m��vx}~`�sn��q������������������||tnjkghophjusoyz{z��z}�~y�}uyus|wu{xx~����������������������~~xuuuqmopoqussvwuwxuuvvtuuuvvwwxz{}}��������������������������|xxvttsqrsssttttutsssssstuvxzz|~���������������������������������~|{ywvvsrrsqrssstuuvwwxxxz{z{}}}~���vw��{���������������������������}|}zywuzvtvvsvwwxuwy~sx�tv�yw|}|w�z}�~{��t��r��x�����������������������~��{x|}wuwxwrr�gv�ze�|j�y{u��p��v}��p��n��x�}�����{�u���������������w��s~�uy��j�{wj�c�ox�X�su�{�d�gu�cz�O��B��p����n�rv�[��b��p���l��k��dt�b��R�gj�ql�ye��o�q�v�j�d�p�U��g�sw�ur�i�ty�w�r�Y��Y��S��i��~~�l��^��i��y��a��e��q��_��[v�M�}ry�[�wi��]�i~�l��mv�M�e�|e�f��s�g���|��t�j���|�p������v��w�z}�c�ue�p�`�o~o�T�ru�sywj�Zr�p�u�k���o�w�m��|y��Z�|�����������j�{a�}kjw`vzml|�gs�ksy�[t��cr�s`~�r`}�rl�~t��q��}����������������|��z{ogokbggfkovj{v~�l�wrw�fxxvllw�`p�~r����||�������������������}rhad\X`V[aijhyxw�����~�~wuyooprsgu}pt��|�}�����{���������������w�~c_YKOVPDN[bcf{�����������}tgh`Za^YX_kpqz����������ŵ�����������|r}p`eRKVVXSUahkmy~�����������xqla`g^Y_\aloot|������������Ú����������{lnoa^MCSWVSSbnu|�����������~wtnfc^\`b^^gkmtw{������������׷����Ʒ�����pkm_Z]A9OSTRZjp������������~pkmg]b_Zbiecmsrz�~�������������ɟ���Ǿ�����xheYS^J:HMS]]fr}���������}|vkfe`ce__fkkoutw���������������է�Ǥ�϶����{wkOO]U>@INZbkmq����������{xvqhh`]ggcfjlouyvz���������������̴�ū�ʵ�����wqYSVYKBKNU_hjn����������~tqrlcadehjijmtxxz}z���������������������������}w`STXULKOQ`mpsw����������}xrmsohjjjrqrnpytz~zy�~�������������������������w�thfabbdfb`iikvuz|�����~{|wwwy|�~}tyomkkmpwz~~���������������������������~xsoifa\[Z[]`fmt|������������~{wsojgeddehjnrv{����������������������������xqjaVNLKLOTZbkt|������������ytpjfca_acfjorvz����������������������������yroh^TOJILRW`fks}������������~xqkheba`_`cglrx{��������������������������{snkg_VOIHJOXainu|�������������{tlfa___`adfjpv|���������������������������~smid_XQLJILT^fnv{�������������|xqjd`]^`behjmrw}���������������������������yojd_\XSPNLNU]epx~������������}ytoje`]]^`dhlqw{����������������������������pfa[YSONOMKQ]kw}�����������~yrnjgcgd\Y_gikpx}~��������������������������}pdZTRRQPSSSW^it�����������zupkhfdccccdfinqv{����������������������������zmaVOKKLOSUW]dmx�����������{vqmifdcceefhilprvz~�������������������ƿ�������zpeXPJHJMRVY]bis~���������zvrmjgeddceegikmptx|�������������������Ǿ�������xndWPJGJKPTX]emw�����������yuqmkigfddddfikpqty|��������������������Ÿ�����wk`UKGDGKOW[`hox����������zwqmjhfffghjjkmmoqruy{�������������������Ƽ�����zkcXLGDFJNYW`fiu����������wvqklgehekkfmkjnqqtw{|������������������п������}wi\QJDBJKQZZbhp|����������zzrkigafkimqkloloutwyy{~�����������������ι�����|pe^LJFELOWabimw�������~xqqppspnrotxvvpfdabinrvux|�����������������ǿ���~mwne`TTW^lnoqa`cbp���||w����zqwqx���zoe^aaenikolq{�������������|�����Ÿ���z�tccPOkhx�ujf]^aihepoz����yjkrt|~x~}~xqd[]_iqywvzy{�����������������̯��yz�yf`X\r��v_YagjrdW[dv����ywpw|zwtry����xg\^bksuysv{x������������������ϭ�yuts{j`gir��{n^VT\abdhq{�����oplgqvt~����{sia`cgqxzwyx{�����������������۴��pottailm���xtXW[]Za^`o�����}rnkrpou|����~{silichllt}xwz~z~��~�����������ɰ�vz�vq`[_w���{aYa^fc[S[q}�����xwxxncmv{����qmhedinpx}}xtyu}����������~����Ԯ�k{�}zmSer���zcXVcgo^]Xg{����xuu~vnjkz����wqplijjktx|z{yvz����������}����׼�~|�}{hWYl��ymZ__jfcUYgv�����qxzzxofns����slihkijjqx|�~yvy���������������མ�~�|v_Sbi~��qhZdeqoe[Zfs�����rv{{{yqmw����sebeirxtquvx}��|{~�������������־��~��z�fVW]gv�|pef]jssmkgir�����yswv{}~{z|yywtmkijlpy{�������������������ʾ����xu�uom]ZZcgnnvmjokot{y~z{vtxvwz|w|z}}�}zzytzzz|������������������������������������zurkjlmmnnnkkonpuvwyyyzz}|}�������~�}~}|||}|~��������������������������������|{vstsrpqonmonprsuwxwxxyy|~���~~~~~�����������������������������������|xwvvussrqqqrtuvwxxxxy{z}}~~}}}|}}}}~~}~�����������������������������������{wvuutttsprrruvxzzz{zz|{|}~~}}}}|}}~~|~~}}~�������������������������������~}uttrrruppptpvuyz~}yz{yy||||~}~}xzx{z��}|~���~���������������������������yvjpknosqrqmqpv~����{vvuw{{{ztxutxy{yyy|y�����������������������������{rpba`adhmkpotw�������}qoloty{ywspnoqsuzwxy~������~�����������������~zwricXTSRZciu{���������������xqniflmrsvqokigloqz~����������������������~ssjd^RONMTbfv}��������||vmnz�~��yrnZgjmvyvlf_]Yll{�����������������©��uxjiZXJJMU^mxz���������}sjdcw�����xmVejqz{te[UQWkp�����������������Ժ���}zree[SMQRUflr|�~������|wmeefu�����|r\okr{uncYSTZko������������������Ƴ��|{uhkaUNNKRalv����������~vommkszz~�zwxuvz{xuoe]^\_px�����������������Ʋ���xwti`[JORXiw{�}tphlrz����vvsv�����yutrvytog\UUXdr�������~����������ƽ����ura\XJRTXeor}yzyv{~�����zuplosw|}~{xyww{vtnd^\]cn{������~��}������׾����|�wl_ZGONWckoqomns�������yohlow~}|tsww|}yoh[WW]ht������������������î��xudi\UUQSZajqs{u}�������|nliiprw{wyxvyvvskga^cis�����������������������~�qj`SPLQV^cifnkr{��������spnnuvyyuuttxwvrjd^\`fr}�����������������˾�����zon_ZUNJQSXchpw����������wpngikkoptstuqppijjjntz�������������������������rqa[SNNRU]adjjrx���������zvvvvxxturppolkgeddinu~�����������������Ⱦ������wvk`ZSLKRQ\ahlty}��������~yspnpopqplmiijjkkopt{�����������������¸�������zrdYPIGIKRZ_iq{�����������yvsomkhgefgilnosswwx}���������������������������wkbWMIIIQV^fot�����������|uqlldc^`^celnwswy�����������������������������sk^XOMKQRY^bnr|�����������~ysngd`bbdfilso|w���������������������������������zqe^WQSTYWb`imv{�����������{xoohmejfjplxp�u�z���������������������������������xpic^[Z^^agcnjyr�}��������vr{mtjsjstvt�w�{��������������������������������ysjifdidj`n`pjxx}��~�v�v�t�t�q�r{vr�p�q�y�����{�l�k�|�������t�u��������������{~qujujtlmpawb{qxy|z}zy||z�y�u�p�v�y�u�s�|������������������~�|�~����������~�~�~�~~~zuzrsuoxnuqrvwx{ww~z{}x�t�y}~~}�z�x�}�}�y�y�x�v�q�z�������|����{�v�y�x�x�w�y�}�x�u�s}xv{u{qq�r�w|}s�p�n�u~}�|�x�s�~~�z��������}�w�p�u�w�{�������{�|�y�z�~|�~|�t�s�{�{�t�l�k�q�u~zx}y�l�e�o�|��|�v�u�{�k�f�l�s�r�o�t��~�~}�v�y��{�q����}�z�{�u�y~�w�y�|�s�k�h�r�r�j�j�o�{t�X�G�=�I�b�~s�a�[�^�_�t��m�u��{�s�u��t�f�g�n�y}�w�~{�x��o�q�}{�w�|v�d�i�~r�q�z}�y�m��z�yv�{|�x��|�y�~��w�s��{���}|�}�����~������xy|z���{yorxx}|ysontw�~zy{w{�z��~�~~���������������~����������������}��}~zw{yvvwsvzxpuwtx|tx}xx{xw}}��{��|������������������������������������}||zyyutwvsuvuwtuywxy{vwyz|{{{|}�}{~��������������������������������������~|{zwvuuututuvvvvwwxxyyzzzz{||}}}~���������������������������������������~|zxwvussrsrsstuvvwxxxyyz{||}}~���������������������������������������}|zxvussqqqqqrsstuvvwxxyz{{|}~����������������������������������������~|zxvtsqpooooopqrstuvwxxyz{||}~��������������������������������������}{xvtrqonmmmmnnopqrstuwxyz{|}~�������������������������������������~{xurpmlkjjjkklmnpqrstuvxyz{|}~�����������������������������������ztokjhfdbbbcfiloqtvwyz{{{{{{{{{{||}~������������������������������wog_XRLHGHLQXair{����������}zwtrommmosx}������������������������yqic\UNHD@@DKS_ly�����������|vpke`\XXY\bjs}����������������������zsnle`YPG?<<@KXgv�������������wl`VNIHKQZdnw������������������������}sk^QG>98<DMWbnv�����������}pf^URPOPQW]dnx��������������ɾ�������}tiVI>8:=HRY`fms}���������{pjf_\VROLQW`my��������������²�������qaL=99@FOVVW\dq���������~yun`UJFIN[gpx{������������²������zh]MFBEGFJMQVas������������qgZPJHPVZbeknx������������ŵ������wdUF@AGJKMPQXi|�����������tdXMJLT^_adfmw�����������ж������cUIEIPQLHKOYm�����������{l[QRSV[]][bmz�����������ζ������y\MPQTZVHAIXfy����������vibZY[ZSSW\ds������������ɷ������u]RW]X[VIFSfu}��}�����ufbcb]ZUOQ_kx������������ų�����zbOP^YZXQKSn}���|x����l[W[\X[XQTiz�����������������tQBLXZc_QL^{����{y����t\LNORU\UTbs����������غ������hHDMU_jbYWo�����|{~}fRIIIQY[U]kx����������¨�����lPIMS`kh`as�����|vwv{vdQFBBMX`_fox���������Ǵ����zgRNOU]beeh|�����~yyuwl`PFCGNY`fjsy��������ȷ�����nYQRWaheefv�����|tssxqaTE@BN^ejnov|������ͺ�����tZOOR^ggfes������ysqvsfXF:<FWcmpot{������ʵ�����tZNMQ_kkkjt~�����wokqng[H=<GVersts�����Ҹ�����}dNGIZiosorx�����riihg]LA;AOarx{y������Ѹ�����{cOBFVeu}~}~������uh_][TNGCGO^n{��������ű���~rcVJKPYht~���������th_TKJFINV\fq�������ʺ����~kYLEHQ]kt}���������uh]RMKIJOR\dy�������������q^MCBGUbmx|��������~o`TPMMRQTWbz������λ�����s_KA=ER^msy}��������o`WPQTUVVbp�������������kXH@BHUbjrv{������vj]VWWWZcky�������������|k[PKGMU[dkqw������wlca_\`hmz��������������xh_WQTTW\bgmv~�����yrkjhghnr{���������������vle\\[\`chkrw|����{vqommnntw}����������������ysnmllmmnoqtwz{{zwtrqqstttvy{~��������������������~}|{z{zyyyxwvutsrqqqrstuvwxy{}������������������������}zxvtsqpoonnnopqstvwyz|~��������������������������~}{zyxwwvvutttttttuvwxyz|}�����������������������������~}|{yxwvvuuttuuuvwxyz|}�����������������������������~}{zxwvutssssstuvwyz|}���������������������������~|{zyxwvuuttttuuvwxy{|~���������������������������~}|{zyxxwwvvvvwwxyyz|}~����������������������������~}||{zzyyxxxxxxxyyzz{|}~���������������������������~}||{zzyxxxxxxxxyzz{|}~����������������������������~}|{{zyxxwwwwwxxxyzz|}~��������������������~���~{wvvwssutpottuvurvwxyz|}�������������������}sokfec_]__]ZZ`ccbdflmx����������������|tfYSPMKNQT^iov���}v}znfa\s�xw��������ŵ�����sic_PGHJMTX\gqtsqw~yuok����������Ŷ������mmm^OKUSSVZdrvqw~wzysmkgw�wy�������Ŷ������|whWQQSHHOZadhozxov~wnkj��tz����������������sfYT^PBJ]YYclsyvj|�ugqn{�us����������������shh^YPGLYTP`mlkrquzskqpo�s����������������zmnaVYKJTXM\jikrupzypothz�su����������������vqt_WWNQTSOegekuqpxuoqne��lx����������������xvt_UZSRPTVdccoupkvyqkni{�mt����������������z�wbW`XPNTX]__orkhwymiqoh�n������������������}kaa]QRUUV__dmkikvpilsfj�xm������������������}idg]OUYTS]`dgghlslinrdk�yl�������������������kjmaPV^UOZd``fkfjnlhoke�m}������������������woqjZU`[NTd^Xbkb`mneiphi�~p�������������������zvri`]`[TXa]Zbg`_mlchslex�vw��������������������|pmkdab_\`b__ed`hlghrrmq~�y����������������������vwxofile^fkbakldhtokrxtp{~||�����������������������~zxuqqqomqroosspqurprtqptustzzy}�������������������������~{yyxvvvussrqooomlmmmmopqsuwy|�������������������������}zywuttsrrqpponnmllmmnoqrtvy{}��������������������������~{zwvtsrqpqqqpqqqqrrrsttuvxxz|}~��������������������������}{yxwvuuutuvvvvwwwwxwwxxxxyyyz{{|~��������������������������~}|{zyxxxwwwwwwwwwwwwvwwwwxxyyz{|}~��������������������������~}|{yyxxwwwwxwxxxxxxxxxxxyyzzz{|}~����������������������������~}||{zzzyyyyyyyyyyyyyyyyzzz{{||}~~�����������������������������~}||{zzyyxxxwwxxxxyyz{|}~�����������������������������~~~}}}}|||||||||||||}}}~~~����������������������������������������������������������������������������������������ao��i|��ty�~|��{|{����z|{~��}����}|�������~���~{�~z�{~�}{��}��~�����w~�vq�z|�v���|�����z��{}��y�z�}�|�~}�}~�|}��~�~~~�~����|�z��{|��{��~~~�}���|��}��|�y~��y��z��{~��u��z}��s��~}���~�|�}z��}}��{���}����~~�}��|~}�|{~�|z�{z|}x�}~~{�}��������������������y{zrnqjfggdgifionmvwv�{���������������������uoke][[UU\ZZ_iihkqxqkx~nmxtz����������þ��������uoiYRRMHHOPP[_dbfqqqpyvqp��~�����¹��ƽ�������p`^VMGIGHMQWcbjlptuuryuio��s�����Ƿ����������}g\TNICCFMNRbghloywruzvek��s�����ɽ���Ʊ����xzd[JKKBCDSUVgmtpq~yvuvoak��r������Ǽ��ǵ����ohdT<BID:CXZ]htus��vosp`k�xy����������µ���xj`XN;@EFBK]bjry�|y��ylmf[t�n~���������λ����obVVB8AIGBWeirx��{{��ndm^Y~xk����������ƻ���wcYRL=<AMLNcow|���}}{j__W]vit����������õ���nZQOD5<HNLXkw}����z�tc_ZPetg{���������Ƚ���~fWFJF:=LYVcs~�����|{wj_ZRFpsX����������ȿ���z\SGII>?Re^g~������xtseSVSA[wlx��������ǽ���}p_R?AGEDMdjr}������|wiZUWK<]xo~��������¸���tg\Q=>GIJTgpz�������wuiZQRO=Vtr���������ķ���udYS??GJOWhq~�������urnXMOPDRrs���������÷���udVQE>ILPZht|�������vqk\QOKFKgt}��������ɼ���yj\RKAHJNZbpw�������xspbUOTJHhr{��������Ⱦ����p_XQDFLNW_ju��������qtlYTPSJUrs���������÷���zk^WMHNKS\cmv�������wqpgZTVQYmq~��������������ueaWHPPPV^ho{}�����|sso_[ZVUest��������ƾ�����ribUQTOSZ^eowy�����vtvkb^^Zcsq��������ƻ�����qlaUXVSVZ_enru���|tvukhda`pwu����������������tsh``][]`bempsyz{|zuvxtqppoq}|�����������������~xuropnoporstvvwvutsrponnpponnpquz�������������������{tmgc`___`bdghiiijkllnprty�������������������wngc_]\]_`bdgjmoonnnnlkllou|������������������~tmhc_]^``abdhkmnmnonlklmpx������������������ypiea]]_abbcfjmonnopnljklqy�������������������vnhc_\]_`aacgknonnoomkjlov|������������������|slga^]_```bfilnmmnnmkjkmsz�������������������vojd_]^``_`dgjllllmmkjjlpw~������������������{rle_]]__^_aegijjklljijlnt|������������������voga]\]\]]_begggijjiijlov~������������������unga]\]\]]`bdfgghiihijkov~������������������woga]\\[\]`bceefggggiklqx�������������������~vmf`][ZZ[]_acddeffffjknt|�������������������|sjd_\ZZZ[^`accdeefghjlqx�������������������zqib^ZXWY[^`bcdeddefhjov}�������������������}umf`]ZYY[]_acceeefghjlrx��������������������}umf`\YXXY\^`bdefgghjmpv|��������������������~vpje`\[Z\^_bdfghiijlnptz���������������������ysnieb`_`acdfhijklnoqtx{}�����������������������|yuromkjihhhhijjklnqtvxz~��������������������������~|yxvutsrrrrrsttuuvvuuvwxxz|||~�������������������������������~|{zyxwvuttttttuvwxy{|}~���������������������������������~~}||{zzyyxxxxxxxyzz{|}~�������������������������~~~}}}|||||||||}}}~~~�����������������������~~~~}}}}}}}}}~~���������������������~�~���]|�h�w���h}�i�zx��`{�{�o�v��f�s�x{�y�t�zy�Z�y��~�~}�{�n�nw�nx�w��j�c��u�t�`�ut�a�i�y�u�c�v}v�P�|p�e�U�vz��w�_��p�|{�o�`�h��f�K�t�v�q��Z�O��uy�m�~�u��z|����u�m��f��{����t�h��v�q�wk�ni�r~Y�Yy�et�k�f�w��[��z�������~������y�{tv�hgqjemafWp{Ltsf~mrz�n��������������������{uykglgf]pahmmkluq`o}cpm|gn�[��������������������}qin`\b]XYe`jfipoclwijqqshm~����������ı������|tnaT^ZUSVZagciojmoski~ieul��}�����������������tlb_WN\RPV^beohqmozfupqkfsk�}��������þ�������upeY[QUUMXX`gljovitsoqokmco�yy��������º�����snkUSULYPSZ_kmplxpqxmtlpn^j��t��������Ȼ������njj\JWMTTR\[npsov{lzvmrkmdf��t��������ž������qffcGNTLQT^[gsutvpt�rhntb]t�w|��������ĸ�����zjcgXBTPMQW^]nuwszn|}ompp_e��n��������ƽ������ufbeOCTYLNb`bsxvvqy�qhsl`l��m��������ƶ������ykfdPERWTLPgektuu|�ru}wvmpjg��s|�������Ĺ�������rmh[PMUYTNWigmruy|~sv~vzqnpm��yx����������������xrucU^XUX\VWnlhpzxt}sw�{~qr�mz�|w�����������������||wjajfZ_eX`qkesypq�uv��vz�|~y{��x���������������������}|wtyuotxtrxvrvxtsusnpqnmqqprtux{~������������������������{xwussrponmkjihfffffhjlnqtw{�������������������������|ywtrqqonnlkkjigggfghiknqrux|��������������������������~{ywtqpponnmlmmlkkkkklmnprsuxz|��������������������������|zxusrrqpppooonmmmlllmmoqrsuxz|~���������������������������}{ywtrrqpppononmlllllmmnprstwy{}���������������������������|yxvtrqqppppoooonnnnnoopqsuvwy{}����������������������������}{ywutrrrrqqqqqqqppppppqrstvwxz|}����������������������������|zxwutsrrrrrrrrrssssttuuvwxyz{{|~������������������������������~}{zywvvuuuttuuuvwwxyyzz{{{||||}}}~~~~������������������������������~}|{zyyyxxxxxxxyyyzzz{{||}}~~~~�����������������������������������~~~}}}}|}|}|}|}|}}~}~~����Nm��[|��^v�{srz�yv���x��z��s��y}�z��zm�s{��l�|~�Y�}�`��f��\�f�f�|x�ll�|~e��i���i�w��hu��rp��qg��S|��pn|�pn��F��y`x��dc��]X��dr��unn��K���fe��uuv�p}�m|��vwx�i|�v���n�{��p{��`��q{��qa��yk���ss��~t���{|{��}����u��{{�w��f���ut���t|��}j�{�xzt}}�}���w���ys�������u������|��}y��zpw�vqbusnknhwpjus|�u���~�����������������������~snvluimmmifquzmxtxy{�zidv|mrnlvrvw�������������������~tonkge`_cehnktpnw�|}yzqhpt}mdfqry||}������������������p`^aaebb_\gnw{ztwz���ufcbktuvsljmv��������������������reWR\bhkhdbgn|���~wyx{|qngkhoplnry}}����������������}uqplf]YUT\emqqrtx����xtpqvniebbm{��}w{���������������}neadfhf_]Z^gty}}yvy���|rmebgnppploqx~����������������~slfda[WX\bekruy~���}|yysoga]]eputqru|����������������ug]WVW\^bcddis|����{vtrnfd`_^afkoty|����������������|l^TOPRW^filnsx����vmc[ZZ\^^_cjry��������Ȼ������p^PHFJQ\isxzxy}�����wl^SNOTZ^cglrwz���������������ydPEAGR^kx�~z|����~uj\PGFMX`finrw{�������ӿ������ygSFDM[iw����yvz~�}uk`SJDIT_fkotz�������������zl[MMTbp|����~wvxvpid_YPKJQ[bflt~���������к��usy�zj[UXan|����|snmljgge_WOLOYckr{���zx������ɫ�tow��vg^[^i|����zogcdjmmjc^ZWSV\gnuw{~wz�����ݿ�tcgv��tkgefs����{kbZYaouqjcb^XTYdknrx��wo������ΨvY[o|�~{woim����~naVQ\q{uokicYTYemmpx�}tfu�����ԩrPSj{����rjp�����q^NQ_s}{xui]VVZ`mv{|zupfs�����̝kLPj~����tms�����nXLRdv��rcYY\afryvqonlfs�����ɘgHPk����xqx����mVP^n{��xm]Y]fdeqxvsrpobm�����˔`EPh|����ww{�����iTXcjv��yf[\`bcm|zolmjga|�����UIUm�����v{|}��}aZbcfv��p``b``jtvphhmlji������wRLWl�����z{tv���veefch|�ugdgaakrmmpojfjoi}�����wLHVl�����zzqs���yidc`ez�vljhcdnpgjqmektpl�����xNHWj�����zwmp��|nha\fy�wokebequkjsmbhsshs�����Ƃ[NO_������xik}���~kfb^kxywskijlomfgmkgp}rf}�����rMENg�����yf`r����rbX\ly~~vldfkrunhlojeoujg�����ݜeKKWw�����tefw����xdca`l{~xqonjmtpbdsnhx{mjw������}XLJd�����{f_l�����f^_]j|�|smjhowzlbhpmqzyoio�����^KMh�����ze[n�����g``[g{�vpmehuyrhipoow{tot�����ݮ}\PXs�����tb`q����zfZ\bmx�uqmjmqttkhotsw{{wut�����ʑl^U`�����}f[i����gY]`gu~ytqlilsroopszzxxzxvx�����Ęyiai������pcky���tb``alz{{wlgimorxxty~wtx{x}������ǧ�ziiz�����zlirx���}oa_`dn{~}{tmjkosv{zty�~wxts~�������ȫ�{hal�����~mmpnx��zth]\doz��skiimy���zwvuw|{z���}�����̲�qb\j�����|gcgmz���xk[[al{���{phgkt~���zuuvvy}~����sv����ձ�p\Vi�����}e_eht���}q_Ycpz���xnkhkw����|rrxvv}�|~��|u����Ͼ�~e\e~�����o`^gr~���zwg`jpr~��}vrkgoz}���{wurpsz�����{nq����Ϫ�kY^s�����s[[ck|���ula_mux��uqmimx����vrmin|�����rpxv{��������yoiy�����tihhlx���~wkiqnp{z{zvnnsw{���~{usqs{�����}yy|��������ª�ygbp�����webfny���yqiemz���~rkpux{~}z{~{zxstz~���yxz�����}|y����¨�l]av�����paair���{tmhhu~���~poros}�{{~~|}~wruz|����}|{y~������{yv}���ø�sa_i�����{g^dmx���woihlu���wtuuvy}~~��~zwtsx����zvz}������~}}������������lhjx�����l[_mx���xljjjv�����uouwz����}|ywz}yz~���}xwyz}����~{|~�����}z}������rcfs�����wh_gs����wkklow���~|yuv{zz�����~|{z|~����~|yxy{���{ww{�����{xwux}������n]\l�����xf_iw���xnlons|����{vssw|�����}|z{|~�����{xz{���|yyz}���|zz}~~|{yvx������cV]p�����sd^n���smonmw����zvvwx~�����~}{wx~�����xsqu����|uuz~������}zyzzyz{zz�����c]j����}rllv~��|wspsvv{�}z{{{}��~|}}}����~}{z}����}zy|�����}xz�����|y{~~}xtsux|�������nku�����yyw{�}utvwwz}wrvxx|��}{{wu|�����~zzyx}�����{z����~��}}~��}{zvux{|}~�������rnt����}xvtz�wvwuu{~vrwxw~�zyzyz����}��|x|�����{xz{|���|~�����{xy{}���|{zvv{�������~yy}�������ywzurx|~|ywrnsyy{~|}~{yz}����|~�~�}{����}uu|����{||zz}~~�����{ts{�������������~z|z|���}|upruuuxyvvzzy{~{x|����}{|�����|zzz~���~}}~{wwz~������|yx{~�������������������xsy}��zxwtuuuty���}vttuuy|����}wrt{����}z|~~~~|}������~}�����|}������������{}������~~}|~}{zyxxy{||}zxvuuxz}~~~|{{z{{z{||}~������������������������������������������������~|{{|}~}{yzz{||{yzz{|}|{{|}}~~~����������������������~~~��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������~�����~yy||y{zz||~~�������������~}}���~~}{{{yz}���������������}||}}~~||~���������������~~~~�����������~~��~~���~~�~~|}~~~�~~~~����������������������������������������������}~~~�����������~~}~�������������~�������~~�~~~��������~~�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������~~~~���������������������������������~}}}{z|}|{{yxyyvvxxxy{|�������������zpoxtjw����~ttsi`gs~������{pkmt|�������{vvxz{~�����|zzyvwz���}}||~��������������������phw����}~�yicjrwyz}���}qnprofgw��|sljkjddoy��|}������պ��xvfZcy�������lWNP[jt|�����vjfdaep�������pc\[Xbw����~wo`VYbk|~��������߸����|UQj����|���fST_lmfk�����}��u]T^p}{oq~��pb`imjfix���������{���������wNRalrysx���ypffk_S[q�������xdZY`lojo{��~sinsllmw��������}���ѹ�����cS]j^^^[y��}|}z�ul]cwyzsuy}}nigmppndjsxumkluuvz{�������������ƾ������|speeaMP^idgliu�vv���tlotoljikrtnou{|~~z}�����������������������������������������~|zxvuttqppvsmnooprrssrtwxy{|||}~����������������������������������������������~|{yxwvuttsrrqqpppqqrstvwxz{}�������������������������������������������������~}|{zyxxwwwvvvvvvvwwxyz{|~��������������������������������������������~~~~}}}||||{{{{{||||}}}}~~~�������������������������������������������������~~~~~~~�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������~�}~~�������������~}|}~{����������~����}~|}~~~}�~~�����~�����|z~�~~�}{~���������������������}~~~~|~}}~�����������������~~�~~~�~~}|}~�����~||{�}|���|}|����������~��{wvy|~���������v~yztw{x��}������������}zvvnqsojmuqtsts��xx��������������{nUZaSA<NN\b\[l����~���jcda`ba_l}�|��������������ȽӬ����xi\LWTH9:OO`Xdq{��������}ttd_NEHKPOUbeu�������������Է���ž�����}_RK>B7,$<OZboy����������thd]K@=@DNONWhw}��������������ž����ѿ�����c[KE>9,'=IPXnv�����������qkeTHFJKMPTVdpwy�����������������������������lTNBH83&4?OR\gy����������vsf[LJMSTST[it{{�����������������������Ǳ�����q`YWK?6<>DIRTbp}�����������~xromnomiinquvyz}����������������������������������xsomligedddeeghjlnpruwxz{||}}~~~��������������������������������������������{wtpmkifdcccccdfgjlnprtvxz|~����������������������������������������������{wsoligecaa``abc