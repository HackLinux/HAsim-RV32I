���b��tK�J��j8����Z���,��DF�i��*��L1�uX�����[	����dw	��,�ęsp��tHY��_zízڔ�k�#s�	_CJ	����D�]*�����gMը�B]����o���*qXU�0y`Pr.ÏY8��&
~�~�����bM�pc�p���P_ԋ��0��*��Е��b �QEaVd0�y>;�
��'E��nft;L�ޚ:��t����Z�q�[�C-e�n�
ك=Q��lǔ<�z��y}�2V\����Qb�Ah
P�+��h^p	M��B�$+�[�_D$\P�+��Cѹݞp,�&��q���+2.�
�B.v��A�F����7�}�rI��+*pT��(K|.�8mb
�ea*��/)��T�g�"|Q�J@��,����@�k  �$aaΩ��$ͷ' �NmFI���`�����{�*��5�Gҹ����31%��e��m$�����7���G
�z�>��S�\n҇&�q�FC��If��Ca_��6�`#7-�����E���\���i��3_�G��G��_-��Iq�ފS�I���$���f��ܮ6y���#�M�`;#�����>k^{řy����?�/�b}"����
"1�@#�DpB���5&컽c�o��!�{I��Úw�"��1���=ߛ���G�W��iڿ������7�^u�_c���b�K�n<�j��~���e����5�q+Q�l�*���^,�G��mb2?2��a���o����Ii�u�L;�ؠ�(N�/�ϟz�/�6��r���06��D�~yM~����e�=x�7P�$�ފ�v"����%���� hJѓQ�qI
�Q�cl�x���a�j��^��=�򎕐GnܧC]��R"���iqg1��YL6��W�Ƴ��W��V���L��V�*�4d�aQ�����?|J#
���6��|<���A���{���	���aڇ_�~A�U��l��t��<k���(��xx��݊�ZEK����5�f���n&��b�+O��:��R�#O_���K�ڰ���\�ʴآ��B��6=�M���#Br��K��ʝ�{R#tq>�g�7b%Z�|�qih�3�l�%��|7�<i��ZRj�9p�:�Ȼn�l-^�/�؊��RĘKju5�h�f��m���!���xs@s�!�,$6��U��&/�5پ��,-��9��
z/�j����،Y�a�Vh7<CK��@�x�+~�t��1ei�[�.b?�J����qV�� �5ǰ������D�Θt����f}��R�؜L[��#��!��~����g�N�۲�P ���&YvX��7����W�$�F�k���22�w�WnǢ���Uw���O��gRs�[���E�cm{ns�W�kK��6�e%�(K�Ǆ�
/��;t�"96y9�kH���)�h!G�"Ř1=lbB[m�W��T�i��E�L[b��։�`�#�g�]c�R�U�`!�gZ�'a��p�ɢd� �MV]�ik��"M'��G-�y�k;��H{KZa�V\/�g|��X�7��ܐ�YVNT,���>�u����zRd7���54U_g�U��2p,A2�9�ͱR��vʃ%�k>�ĖF�X�H��T��x�b<�?�U6�y��i����QV��$|T&��I�3�N/�<d̢E3���i˕����3X�j���ҀwFt��v��d�8<��;(�I�ꎕ��F?Y���\���)3��bI1N�9�]����>7$���&�P����>�>�i�T�J�q}��h声�H��aQ�qz�&�:5���م��Q��kIQVNr�E�M�D�)���-�ʈ�eLa�E-�׻>#��lӭ�ף,�8���U8��S"�
�-7'�0��{������k��h�?��3T_K�F.R���Φ�J�+��~�Ϗ�F��OخVsm�<�ڻb��lau��su������}���̒@�y	#)��W�a�y�J��IR�g�x������D�41���@�,(�|-Ĵ��V�ن�fi�G[f�i����aX�\2���'�i�o�l�Z���	ț/H�4���;�-W�c'�������`/���Y+ʐ�s)O壐9@� A$�x����3{�hw�7X����&[���".Xٛ�M�ѕ�AWC�=s�{��z���eJ`�R�csQtjWU�;{@@�ŹQY��n���Ёn	m킥ܼ���-4�8ID�VHc˫�l���T�����S�b,$�u���6=]{��Wj]طQw�E�X�~�Ӡ+&սA����@���=�	���hmpw��=v�Qr�ՠ�ؗ��N�2��(��{�L�<{h�?y�D���qQK�>�(�[hԼˏ�����yZB�V���h �4��S��)AU�D�2�Xw3튴�M󓤎o�cպ�_�'��x�	��n/�9�;+�/l��C%n|�E�#��5\Hob�U]{���t����遝�!R0����_��ǒ}�Q�M-멉.�Q]�:˯��\��'�B�96����̟T���B�WuF��1A��NC��i��`�^���C-�];�Y7�^�����@��Z{)�Q�M)��A��ñ�[�g�Ha�^���i���+F���Z{�#v����#�zi�6�����9���2��C�g��ݗa<�J�.�'��-c�g�ɞ���������ac�Q�v��
%�6��{���	i��eF��c����F�N����<^+Y�Yi/���R5�d���=������7�9�O���"W��'��f�tI1���Ĥd�
eE/%֦}T�ZK��6O��9�!��.rM�t���^v`elS�X47�?Z�;��<���oC��0/@c��$��K
� �1g�ދ�t�jv/M�aQm�̆qt53ޔu˲)������7߰}��W[0�-��|���/�g���bb�g���~4�<�[(ب� �J��A/�pv�k#Ky��4�*8yD��|���IT��nvF����x��6ػ�T�_h���F��9:��v�S)�8C�vs��n�2zK�o͎�ÈB�Br��"�oE�|e��O�2��h�� ��hJ�­�(�hKӹ<��P�AY�͸�vo.?Kj�]��	ue�(��\���QI���1
<w{~�o?���G;�i4����T[�r�u|�n���:���R��f�cs��7��חC;�����h���	V��QN�2ᇊ���I�J���ϭ���Je�S[��8�ۦ�0{W�`�Q��HF�����	SQ��kyS��Q�^Į�r��5�:�]JG��,�7O �z���թ��H��-��l|"-T�5�ut�0�R��	�xn�����,�Ѣ��ʇ4��
W�a��y��Hp	���/��=�0��t������Z�����#U0Z��;���;�rْ�'�l����!�}�F[�5Eߗj��^�;FB���IPd�.��qN���!P��!��n���1
I���6���v)�).��,TZ�<�)0�?�����:�MK���3�<@�!�� A��O|!p"����G9ʦ�-�1��h���e�� ib�}Y�ʾ2t�ῄ��L���Ax���Rڰ��bX�PM���KRtFY�hi����+�דvb1�M���t<�-Rxc�_ye=d�:������~B�����8�!Z-���D�44v�!���*�p;sw�,���;	ZPG�vv�z�[כ�������W�>�`��	$�61���D+���0��uX�6�f��{ڔ.���'���ȢCL@��+V43M�XWt�YW���*J���1��\�"�����86@�tŝ.�!�3W&6ŹP�1|]�~�̊����۳���v���4�Abjzns� �;#g�6�9o�j�WW��)�JL�b���635�����i�P��䝵��a�μņ���0�*���JW���6�4�kS����˟��i�*�[2-0�I����j���-Z�U���T�O������7�o�����ʹ��.�68���� �,;Yr$9�	 dim��VJl���J�Ekh9J-%���(��@K
�����҃�@����7