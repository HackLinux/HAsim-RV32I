Q���]� ������U���(�M؋E؃x ��   �M؋Q�U�E؋H�M�U�U��E�E�M��M��U��U��E�E��	�M��8�M�U�;U�t�M�����3�����t�M�Q艇
 ���ЋU؋E؋J+H����8   ���E��U؋B�E܋M�Q�Y�
 ���U��B    �E��@    �M��A    ��]���������U���L�M��E��H�Q�U�E��H�M��E��U��B��u;�M�M��U�E�
;H��ڈU��E���t
�M��U��	�E�H�M��U��U�뺸   ��t:�E��MQ�U�R�E�P�M�Q�M��s;  �E̋Ű�M��U�E�B�E��   �M��M��U���u�f�E��H�MȋUȋ�EċMĉM�U�+U����B��t5�E��MQ�U�Rj�E�P�M��;  �E��M���E��M�U�Q�E�m�M��� �E��M�P;����ȅ�t7�E��UR�E�P�M�Q�U�R�M��:  �E��E���U�
�E�MۈH�E��E� �U��E��M�UӈQ�E��]� ����U���<�MċEċH�M�U��E�M�M��U+U����B��tG�MċQ�U�E�E��M+M����A�х�t&�M���8  �EċH�M؋U؋�EԋM�Uԉ�E�K�E+E���@�����A�х�t&�E�EЍM�O  �MЉM�U�R�E�P�M��ɻ ���M�U��E��]� ������U����M�E�H���M��U�BP�M�Q�BP�M��8  �M���U�B�E��M�U��Q�E�H�Q�B��ug�M�Q�B�E�M��B��u
�M��U���E�H�M��U��E��M�Q�B�E�M�Q�B��u�M�Q�U���E�H�U�Q�#�E�H�M�U�E�H�
�U�B�M�Q�P��]� ����������U����M�E��M��U�E��H�
�U��B�H��u�U��B�M�H�U��E�H�J�U�B�M;Hu�U�B�M��H�-�U�B�M;Hu�U�B�M��H��U�B�E��M��U���E��M�H�U�E��B��]� �������������U���P�M��E��H�M��U��U��E��H�M�U��E�M�M��U�R�E�P�M�Q�M��M����U��B�E��M��Q�U��E�P�΂
 ���M��A    �U��B    ��]��������U����M�E��Q��t�q�E��Q�B��u,�M��B�E��M���B��u
�M���U���E�M���5�U��H�M��U��B��u�M�U��;Bu
�M�U���ӋE�M����]����U���`�M��E��H�Q�U�E��H�M��E��U��BQ��uB�M�M��U��R�M�^p��3Ʌ����M��U���t
�E��M��	�U�B�E��M��M��3҅�t:�E��EP�M�Q�U�R�E�P�M��;  �EȋMȋ�E��M�U�Q�E��   �E��E��M���u�f�U��B�EċMċ�U��E��E�M�+M����A�х�t5�E��EP�M�Qj�U�R�M��;  �E��E���U�
�E�M�H�E�z�M��ˋ  �U����U��EP�M��fo��3Ʌ����х�t7�E��EP�M�Q�U�R�E�P�M��:  �E��M���E��M�UۈQ�E��E� �E��M��U�EӈB�E��]� ���U���P�M��E��H�M��U��U��E��H�M�U��E�M�M��U�R�E�P�M�Q�M���8  �U��B�E��M��Q�U��E�P��
 ���M��A    �U��B    ��]��������U����M�E��QQ��t�q�E��Q�BQ��u,�M��B�E��M���BQ��u
�M���U���E�M���5�U��H�M��U��BQ��u�M�U��;Bu
�M�U���ӋE�M����]����U���,�M܋E܃x u	�E�    ��M܋U܋A+B��8   ���E؃}� u	�E�    � �U܋B�E�M�M��E+E���8   ���EԋUԉU��EPjQ�e�M�U��M��<  �E܋H�M�U�U��E�k�8�M�ȉM��U�E���E��]� �U���,�M܋E܃x u	�E�    ��M܋U܋A+B��T   ���E؃}� u	�E�    � �U܋B�E�M�M��E+E���T   ���EԋUԉU��EPjQ�e�M�U��M��oE  �E܋H�M�U�U��E�k�T�M�ȉM��U�E���E��]� �U����M��E��@    �M��A    �U��B    �} u2��c�E��0�}� v�E��E���E�   �M�;Ms
�M�����3�Uk�TR�ч	 ���M��A�U��E��H�J�Uk�T�E�P�M��Q���]� ������U���(�M؋E؃x ��   �M؋Q�U�E؋H�M�U�U��E�E�M��M��U��U��E�E��	�M��T�M�U�;U�t�M������3�����t�M�Q��|
 ���ЋU؋E؋J+H����T   ���E��U؋B�E܋M�Q��|
 ���U��B    �E��@    �M��A    ��]���������U����M�E��M�U�E��M��?N  �E��]� ������U���d�M��E��H�Q�U�E��H�M��E��U��B%��u_�M�M��U���UċM�,o���E��M̋M��o���Uċ�EȋM�;M���ڈU��E���t
�M��U��	�E�H�M��U��U��3���t:�E��MQ�U�R�E�P�M�Q�M���M  �E��U���M��U�E�B�E�  �M��M��U���u�i�E��H�M��U���E��M��M�U�+U����B��t8�E��MQ�U�Rj�E�P�M��M  �E��M���E��M�U�Q�E�   �M��+�  �E����E��M��n���M���U��M�
n���E��M��U�;U�����ȅ�t7�E��UR�E�P�M�Q�U�R�M��M  �E��E���U�
�E�MۈH�E��E� �U��E��M�UӈQ�E��]� ������������U���P�M��E��H�M��U��U��E��H�M�U��E�M�M��U�R�E�P�M�Q�M��=K  �U��B�E��M��Q�U��E�P�.z
 ���M��A    �U��B    ��]��������U���(�M؋M��?Q  ��]������������U���,�M܋E܃x u	�E�    ��M܋U܋A+B��4   ���E؃}� u	�E�    � �U܋B�E�M�M��E+E���4   ���EԋUԉU��EPjQ�e�M�U��M��Q  �E܋H�M�U�U��E�k�4�M�ȉM��U�E���E��]� �U����M�E��Q%��t�q�E��Q�B%��u,�M��B�E��M���B%��u
�M���U���E�M���5�U��H�M��U��B%��u�M�U��;Bu
�M�U���ӋE�M����]����U����M�E��M�U�E��M��[  �E��]� ������U���d�M��E��H�Q�U�E��H�M��E��U��B!��u_�M�M��U���UċM�<k���E��M̋M��,k���Uċ�EȋM�;M���ڈU��E���t
�M��U��	�E�H�M��U��U��3���t:�E��MQ�U�R�E�P�M�Q�M���Z  �E��U���M��U�E�B�E�  �M��M��U���u�i�E��H�M��U���E��M��M�U�+U����B��t8�E��MQ�U�Rj�E�P�M��aZ  �E��M���E��M�U�Q�E�   �M����  �E����E��M��*j���M���U��M�j���E��M��U�;U�����ȅ�t7�E��UR�E�P�M�Q�U�R�M���Y  �E��E���U�
�E�MۈH�E��E� �U��E��M�UӈQ�E��]� ������������U���P�M��E��H�M��U��U��E��H�M�U��E�M�M��U�R�E�P�M�Q�M��X  �U��B�E��M��Q�U��E�P�>v
 ���M��A    �U��B    ��]��������U��j�h�-' d�    Pd�%    Q�M��E�� �p( �E�    �E������M���'( �M�d�    ��]�������U��j�h�z' d�    Pd�%    ��P  ��?3 3E�E艍�����E������E�H��`�����`����� @  ���G  �E�P�M�����������������������E�    ������R��������E��E������M�����j �M��� j j�M��~x���E�   �E�P�M��������������������,����E�j�j ��,���R�M������E�j�M��T� j j�M��H'����h���P�M��������������������(����E�j�j ��(���R�M��`����E�j��h������ �}�r�EЉ������	�MЉ�����������Rj�EP�MQ诚  ���E��E�����j�M��� �   蹟
 �     ��d���R�M�I����������������������E�   �M�Q������������P������Q�UR�EP�M�Q�%Z  ��P�U�R�E�P�
�
 ���E��E�������d���������M��U�;�t�(�
 �8 u�}�w�E��E��MQ�M萨  �Ѕ�t�E ����U �
�}� }�E ����U �
�3��}� ���M$��U�E��M�J�E�M�d�    �M�3M�ͼ
 ��]�  �������������U��j�h�z' d�    Pd�%    ���   ��?3 3E�E���(����g�
 �     �E�P�M�������$�����$����� ����E�    �U�B�E��� ���Q�U�R�EP�MQ�U�R��X  ���E��E������M�������EЃ�-u�Mщ�����	�UЉ����������E̋M�Q�U�R�E�P膝
 ���EčMQ�M�>�  �Ѕ�t�E ����U �
�E�;E�t蘝
 �8 u	�}���  v�M ����E ��,�MЃ�-u3�+Uĉ�����	�Eĉ�����M$f�����f��E�M��U�P�E�M�d�    �M�3M�H�
 ��]�  ��������U��j�h�z' d�    Pd�%    ���   ��?3 3E�E���(�����
 �     �E�P�M�z�����$�����$����� ����E�    �U�B�E��� ���Q�U�R�EP�MQ�U�R�\W  ���E��E������M��G����EЃ�-u�Mщ�����	�UЉ����������E̋M�Q�U�R�E�P��
 ���EčMQ�M辥  �Ѕ�t�E ����U �
�E�;E�t��
 �8 u�}��v�M ����E ��*�MЃ�-u3�+Uĉ�����	�Eĉ�����M$�������E�M��U�P�E�M�d�    �M�3M�͹
 ��]�  �������������U��j�h�z' d�    Pd�%    ���   ��?3 3E�E���0����g�
 �     �E�P�M�������,�����,�����(����E�    �U�B�E���(���Q�U�R�EP�MQ�U�R��U  ��P�E�P�M�Q誚
 ���E��E������M������UR�M�j�  ����t�M ����E ��M̍U�;�t
�
 �8 t�E ����U �
��E$�Mȉ�U�E��M�J�E�M�d�    �M�3M蟸
 ��]�  ���������������U��j�h�z' d�    Pd�%    ���   ��?3 3E�E���0����7�
 �     �E�P�M�������,�����,�����(����E�    �U�B�E���(���Q�U�R�EP�MQ�U�R�T  ��P�E�P�M�Q葙
 ���E��E������M������UR�M�:�  ����t�M ����E ��M̍U�;�t
蒙
 �8 t�E ����U �
��E$�Mȉ�U�E��M�J�E�M�d�    �M�3M�o�
 ��]�  ���������������U��j�hhz' d�    Pd�%    ���   ��?3 3E�E���,�����
 �     �E�P�M������(�����(�����$����E�    �U�B�E���$���Q�U�R�EP�MQ�U�R�|S  ��P�E�P�M�Q苛
 ���EĉU��E������M��S����UR�M��  ����t�M ����E ��M̍U�;�t
�_�
 �8 t�E ����U �
��E$�Mĉ�UȉP�E�M��U�P�E�M�d�    �M�3M�6�
 ��]�  ������U��j�hhz' d�    Pd�%    ���   ��?3 3E�E���,����ח
 �     �E�P�M�j�����(�����(�����$����E�    �U�B�E���$���Q�U�R�EP�MQ�U�R�LR  ��P�E�P�M�Q�r�
 ���EĉU��E������M��#����UR�M�נ  ����t�M ����E ��M̍U�;�t
�/�
 �8 t�E ����U �
��E$�Mĉ�UȉP�E�M��U�P�E�M�d�    �M�3M��
 ��]�  ������U��j�hhg' d�    Pd�%    ��   ��?3 3E�E���h���觖
 �     �E�P�M�:�����d�����d�����`����E�    ��`���R�EP�MQ�U�R�	W  ��P�E�P�M�Q�Q�	 ���]��E������M������UR�M跟  ����t�M ����E ��M��U�;�t
��
 �8 t�E ����U �
��E$�M���U�E��M�J�E�M�d�    �M�3M��
 ��]�  ������������U��j�hHg' d�    Pd�%    ��   ��?3 3E�E���`���臕
 �     �E�P�M������\�����\�����X����E�    ��X���R�EP�MQ�U�R��U  ��P�E�P�M�Q���	 ���]��E������M�������UR�M藞  ����t�M ����E ��M��U�;�t
��
 �8 t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    �M�3M�Ʋ
 ��]�  ������U��j�hHg' d�    Pd�%    ��   ��?3 3E�E���`����g�
 �     �E�P�M�������\�����\�����X����E�    ��X���R�EP�MQ�U�R��T  ��P�E�P�M�Q��	 ���]��E������M�������UR�M�w�  ����t�M ����E ��M��U�;�t
�ϓ
 �8 t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    �M�3M覱
 ��]�  ������U��j�h�z' d�    Pd�%    ���   ��?3 3E�E���,����G�
 �     �E�P�M�������(�����(�����$����E�    ��$���Rh   �EP�MQ�U�R��M  ���E��E������M������   ��t$�M�Q�U�R�E�P苒
 ��3ɉ������ ���� �U�R�E�P�M�Q訕
 ��������� ���������Uċ� ����EȍMQ�M��  �Ѕ�t�E ����U �
�E̍M�;�t
�\�
 �8 t�U ����M ���UċE$��M�U��E�A�E�M�d�    �M�3M�9�
 ��]�  ���������U��j�h��' d�    Pd�%    ��<�M�j �M��س �, Pj �MQ�M��|���E�    �U����U��E��P�M��  �E��E��E������E��M�d�    ��]� ���U��Q�M��M�������E����t�M�Q��e
 ���E���]� ��U��j�h��' d�    Pd�%    Q�M��EP�M���  �E�    �E������E��M�d�    ��]� �������U���<�MċEċH�M�U��E�M�M��U+U����B��tG�MċQ�U�E�E��M+M����A�х�t&�M��e^  �EċH�M؋U؋�EԋM�Uԉ�E�K�E+E���@�����A�х�t&�E�EЍM��I �MЉM�U�R�E�P�M��yX  ���M�U��E��]� ������U��j�h��' d�    Pd�%    ��   ��X����E�$I��}� v�E���T����
ǅT���   ��T�������X���;JwUj �M��̱ h�, �g
 ��Ph�, �M�葒���E�    �E�P�M���m���E��E�X/( �E� hT�- �M�Q�	�
 j �UR��X����HQ�UR��X����HQ��X�����]  �E���X����B����X����A��X����E;Bu4��X����Q�E��B��X����Q�U��E��M����X����B�M��H�e�U��t4�E�M����X����B�E��M��U;u��X����H�M��U��E���)�M�U��Q��X����H�U;Qu��X����H�U��Q�E��E�M�Q�BD���m  �M�Q�B�E��M�U��A;��   �M�Q�B�H�M�U�BD��u,�M�Q�BD�E�@D�M�Q�B�@D �M�Q�B�E��R�M�Q�E�;Bu�M�Q�U�E�P��X����E �M�Q�BD�E�H�Q�BD �E�H�QR��X����F �   �E�H�Q��t�����t�����M�U�BD��u,�M�Q�BD�E�@D�M�Q�B�@D �M�Q�B�E��]�M�Q��p�����p����M�;u�U�B�E�M�Q��X����E �U�B�@D�M�Q�B�@D �M�Q�BP��X����D ������X����Q�B�@D�M�U���E�M�d�    ��]� ���������U����M�E�H�Q�U��E�H�M��U��BE��u8�MQ�M����O��3҅�����t�M��Q�U���E��E��M���U�뽋E���]� ������U��j�h�' d�    Pd�%    ���   �� ����E�HU��tUj �M��7� hL	, ��c
 ��PhL	, �M�������E�    �U�R�M��Yj���E��E�@p( �E� h�- �E�P�t�
 �M�M��U��U�M��}  �E��QU��t�E�H�M��'�U�B�HU��t
�U��E���M�M�U�B�E�M�;M��+  �U��B�E�M��QU��u	�E�M�H�� ����B�H;M�u�� ����B�M�H��U�;E�u
�M�U��	�E�M�H�� ����B�E��M��;U�uS�E��HU��t�U䉕����&�E�E��M���BU��u
�M���U���E�������� ����Q�U��E��������� ����B�H;M�uP�U��BU��t�M䉍����(�U�U��E��H�QU��u�E��H�M���U�������� ����H������Q�	  �E���U�Q�E�M����E��M�;Hu�U�U��=�E�H�M�U��BU��u	�M�U�Q�E�M��U�E��H�J�U��B�M�H�� ����B�H;M�u�� ����B�M�H�2�U��B�E��M��;U�u�E��H�M��U��E���M��Q�E�B�M�U��B�A�M���T��x����U��T��t�����t�����������t�����x�����
��x����������M��QT���  �	�E�H�M䋕 ����B�M�;H��  �U��BT����  �M�U�;��   �E�H�M�U��BT��u&�M��AT�U��BT �E�P�� ����X  �M�Q�U�E��HU��t�U�U��   �E��QT��u�E�H�QT��u�E��@T �M�M��h�U�B�HT��u(�U��@T�M��AT �U�R�� �����X  �E�H�M�U�E�HT�JT�U��BT�E�H�AT�U�R�� ����X  ��   ��   �E��M�U��BT��u%�M��AT�U��BT �E�P�� ����X  �M��U�E��HU��t�U�U��   �E�H�QT��u�E��QT��u�E�