 �   ���������������������  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������  ��  ��  ��  ��  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������  ��  ��  ��  ��  ��  ��  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������  ��  ��  ��  ��  ��  ��  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������  ��  ��  ��  ��  ��  ��  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������  ��  ��  ��  ��  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������  ��  ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������@@��@@����������������������{{��ff��bb��{{��������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������))��  ������  ��CC����������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������������������xx��  ��44������������

����������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������������������������������22��  ��������������^^��  ��xx������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������������������������������������������  ��MM������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������������������������������������������  ��..������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������������������������������������++��������������������..������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������������������������������������������������..������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���������  ��JJ������������������������������������������  ��..������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������  ��..������������������88��  ��������������^^��  ��BB������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �������������**��  ������������������ii��  ��QQ����������**��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   �����������������??������������������������������  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ����    �������������������,,����������������������((������00����������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ���    ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���� ��� ���    �   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   �   ���� ��� ��� ��� ��� ���    �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ���� ��� ��� ���         TRUEVISION-XFILE.                                                                                                        