d��fNU�²�e ��q3+M��جr�,w���KN��m���ɖj��5kv��'r��4���Qψ�y*I��2R:�O�Y��H�)��;�8UH��.�e��zR��0E�g[�BybKA��E,�h�<�$�k� ljZ-vד�e��c�~�e4Y�le�F-M�yIu6;��V��e�#M�L�P)����b�o�n���Q74���M�ў��pT�|FҢ�r(;���������j���8��n畡7h)��6�$�����cs�*v���iI
�ZbQ��"Ka��nZ있�m7��E���q�AH�r�n�,"�Q*�&9����g��{�4������<��O�AA�s81�޳���O��Z*_�r��_]-KάNnn7�a�,��m���:�W�@�Ac�j����8�U'M[M�jW=���߱��,�yj��7}�@�P�7����Q�;b�nx^�Lk�F�F��R�[�X2nz	se�Ĝ�L\���C���u��)�LoڰQ�ц��X�R�+�ʄ䤮p1ٺb�ݮ����@���X3K)2�	얱�~Nv�w1<:2ʆU�2�1��JW1(©$���J�=1A��37����O@��Q��^Z���xuO��)Oz��>����T�j�3�<Z�-�1��9m�����ZjD��z�#��,�u���ps5��o��L��=g�X�..����j�k*yO�WQ/�|/�#�'FC�j=��z��ݹɩρ\ %�Y��G��h_�[����d���7�,Yٳ�
J~w�޵���ו)��D7EjED�7h4�h��:��680ޔWl���5���F̽��Lk��i�!aހ�Mwt���ˀ:yb͢Q�'~�l{�mR��=�Vk�f��eV���Lϥ]�Vl����,��ٝ�fV<i���`�y�U�o�0����v0oN��1��J	#Aʹ��i�Z1:�"O���>��v�\���्%7��#1�UǢ�QM�A�a�/N��,��n��)R5�Fz��� U���h�0�����L���̅&��5ǩn]�_D[KT@GY.�ʳr���C�kh�]-9��uJ���2��X}]�j�-��c���`����s�*|�.��ٿh��|u�25�X�}�m�s<�k\���]�R>���;y�F�e%��7���\(��ң��JH�z.,VR*�&�Q��o���&8���x�T6LU��N{�	H2붵�'sNFx\'-��u9�Z��g��N�N�͜ղs*��m�hK7Q�%���ǖ$�]���]WM%��S�9�c�Ef��%��f,�4��uAOչ	����#Н�5qR#�b���Uӷl��*24n�w������)W[��8�\�V�^�r��ل�]N�v*�xm؄�^���r<�sS/�W�O%7�b���[E���J��l�	�E��@n��%ٸ��Q�۵v��2���2/k8����u����H3�˲��t�]�z�c���0ج.���h��b��Z�tY��%�\�d��+g��dX�,�$���ʩ�rSmNα��6�L���)�Hc[�|��PN�u�w_'Z�ʲNt����{+�ip�R��/�:?��O��U��̦���#�
8aW�T�Q%�zv~z��1��t=�ՏJ��{�����b��ߏ_Y�ak3���͙������q3�������q�����_�י7�2{��mU�DgX��P��ب��G�(}f�GU㖨�єa��&|��	�q�5�1���{�u�މw��޾��̈�NU	Kzi������l�^����������]{�������B/'�{��^�ҡr�q�> 8 �  1`$  Y +%D�?�GRWy�Zz�U>Iw��uwu�np�D�B���,�PC"�l/k��2fV��h� ��@�  ���JS#�@�j���8��5�U�Tl�]��V�2��=�jl���e�Z�M󴕬֪�k̥-��,�t: �w �  H �f� ���ֶf[!2Q"\���*��#������<�$p�-�XHHʫ1WB{ ���o-'��C��>p���鑇�h@�@\����*2��� �0P�/}u��"�U��`@���V%oG5Hr� ��8k����i�8��<��/�F/�ց�Z��D�O�u�LHϡ�
�p)kEp1 �C��Y���8w-m;k�b<|L9~� ��#$�E����^�u�S���AuBn%]_�Yu���k�;$�5 i��KU��0���8����JkBr��x1���C�h����`ʀj�`5�ʇ@��G'�E�~�r���(�ߞ��y��Ň2����8�2d�B�}��T$�'D��a�Х����}l��`����^H�&�[�2JP,9?��|���2����b�]��cb�҆�!����W8|�7��{�`U��*0g�z���E��B�{�ٓ������g�Ik�99���[?
U�#J�9I����,jk�}�q��������r��s5V|A��Aj_�ve�qѱ��s��$�`w3��� �=���v�%}����d6�ᝌ,x�\�����7o���V�u�㋽!7���@����r�w��ǍL
�o�߉��(td�N��YOt��]�kO߯�_m����<��TۋP�
�J"�{�m}� 럢�2��=I֋V��T_�cQ�;ac�bHف��>=Lm���孴�~���6di�� �Jwtl�C�4�W�J�x?8_|!9�t����b��?���o��p�{V
!!+�R�'���}�/�X��<$�:"g��\y�ܱ*lPe=�Jm�j�����7*����@B��x2�)��Tߕ_@|�O�x}��(��-��lރUq$�%
�wE�#���;	�}����!�����\D{P�qD|v�|"}
��f�Dt�$/,�#$��P��V�SVW4�z���8�8��,�=y(�x�@�=#���y�KQM������<�K;IO'�,&R))�4I�����������K�F��/n(�B16��F=��3e�:�*��W$��+cڏUI<:�Wb��͏�s��
�������q؀	��Z���Eq4tL�b����7:�E.�ȅ�؏���ӆ�Q��\��ׯ�SH��6��������,��>��f��@�� @�'|aV�������X�*Y���ӥ�x_����mO+��|����9���.Rw�QOt��M��DݏO�&Gu�����E�@�Z$�)P�&�U^��/�����QF�Ԑ{{�x@���v.)��w�HCn\������{X@[@4h�3 �o��8��_G��|�@@b���{_3Y�� *HH.
}�aZ.7	��
�	b�E��@j�xO��Z�'{��K~�{ÝIA"db�~d«��\������w���� UC�}������AT�C���ȵ$ϑ[��6�ޕ�J��D�� 7��y��%���#�~~�x�g�*��l?gK_u$?��P���8d-wR���
��y�$��|�w��~����]�t�Ewr� ����i��},;��
�{E$�	�Â�u�����mn��si���xܴp��,���O�{��l��D���Eb�*P�~�ߍ(�p�������y�N�|? 9kv�l�C���_�}b�NW ��0����A��}d�}�!K�����V��'
���Ɵ���m�x�x��e�$�{`/$�`yP�3��oy���*�x9�B�"�7���/��\��N��+^܄7���7 7^g�z�㬰���,%�N���o�xp[xC6�d��X���c�!�.: �t�;
̄�@�2�de�,�*��H4y��)�՗A�V�_$O�O�?�Q˺��I�#�G��B����`ܳ�'��á*��˷	F�������v������rmp���Ӏ-;�&�S}�0k�$�=����i|\�7�ȧzg��!������`K�����cf�m`�K!LRP*�����/�н?�y]X	h�Ũ���c¸{R��ֿ@"��J�����_HD?��ل��/2/]A_P�0q��d�7��>9�L�J�_��l%����1��0�XdϝU�Z*_r�<�.ms����PP��e|}��(�H0� G�|����pXv��t?*7�[��j��?>J���Ŕn4�JM����ǚ2�X6z�f8�$yGd�_@y�Q"G��= �ŰӼ=�����y̓����J	�4��X����"���������X�*�O�#����vy7zg