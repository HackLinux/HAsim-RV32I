��(���u�
n	o	�
ER��
�	/6o/��Dw�|�C	z, <$�#))q�����!#P&],'''U())M(�$�$+&�'�'^&�'7)�)�)�*�+>-�+�*`,�.j0�/�-�'��!F-6�0))��^���-�<�����A�����"ԕ�o�����́�ɇ�Fϱ����(�a��]�+�w����ö��͞�0ِ�����))��@�ǳL�d�0����ո��՞:����H�`�O�U����޻��b��]Ǟ��D�Җ���'�m�T���E������9�$~�
  �
�
�
$��D�% � n  ��>���6���"���$�"�Y�����w��C���%�j� ))\ T�D����0D���>����Հ�@��b�������Z%�*�.�0� �:Y"�-8]�C�����Tk))s5�z��2������:�+�pe� ��
��n�@ݟ����{�����\�=��9��:G'��))d���tZ����m�O�S�����U�	IX���& �������<���}�?�G��<���<��I�p�   �                  t�*          �      �J�      t�          8      ��X          �                    l      ���	     	x	�	      
�
�
          H      ��P    T�      P�           |      �N      ��X            33  ��� � � � z n b S D 4 $   ����������������������������������������������������������������������� 	� � � � � � � � � ##� � � � � � � | p g ^ U L B 9 L ^ p � � � � � � � � !#�  ����    	          ����������������������������          33��������~&�E�d��R� � g ?    ��������������u�j�a�X�P�I�B�<�7�2�-�)�%�!���������	�3!@( % # $ % % & ' ( * , . 1 4 7 ; > 9 4 / * & "               2�.�,�1�2�1�0�.�,�*�(�&�%�$�##%�(�+�/�3�@�P�_�l�w���������������j�T�?�*���������������������������33	�������d����f���=�}�����������������{���	���e�	�������;�������\���9��H���w����Z���������K�����33p ����X��� � �Cl���4��-?�n��+�g��������������[����j�J�9�6�<�G�Q�Q�;����������P�33:�5�1�M�N�M�L�K�J�H�G�E�D�B�A�@�?�>�>�?�?�B�F�J�N�Q�T�W�Z�]�_�X�P�I�B�<�6�1�,�(�$� ���������"�33����������������������S)����lP��<u��N���!7<0��33���5 ���/�o����V���������Q���t�������������'���S Z y n @ ����+���&�����e���?���e�)���������.0����������������������������������������������������������  ������������������������������������33������������������������ +7DN8"������xfUE90.2<IY33t���<������w�������7���(�����8�����9����������T�������_��Q��&��Z�����U�#�������D�����.���X���33��l�9�g���� U"� �������:�{���-����d�����\�������h�P��a�h����A������x�Z�=�����[���v���n���$j����� � �"�'�-�3�9�?�D�H�L�O�R�T�V�X�Y�[�[�\�]�^�_�`�a�a�b�c�c�d�e�g�h�i�k�l�m�n�m�l�33������������������������������������������x�:�������s�J� ������n����^�����D������N�������������m�3�33��	)���\"$4:3���oK:H�RV����h	�	�	�	�	�	m		�[�|�&�f"����y33  �]�3
(�		z�8�	}�s�i�D��  �����d�8�8�q�����������L���&���"���$��������8�~��� �<�u�33  ��������z�����z�G����F �i��	�
K�T\&����k�2p����9`
�	�#��5��33  � �](�����0 �_�g
�6f�������!�#J%�&�'\(�(�(�((h'�&�%�$�#�"`!( ��J��$����3��3E�( �(�f�
b�V�&�u�)�'�U����z�5�x��Ω��ώ�p֯�Y�X�A�
���-�r\�M�d���,�3 (������
ջ��9�qҨ��б�Z�
�,�4��%҇�X���c����0�>�%�(�(�(�(�(�(�&�#! ��( ����P�I`�I�/u��/�
�
+
�� I-�������� ���	�	�	�	�	�	��� Z�(� '5�Yp&p �"3&p)z,S/2�4�7�:�<	<X;W:9*7^408)��� �m�Z�B���e��֯���z��l������b�33C���	��TdS_��  a!����	��l���!�g�����W�=�e�������-�_�����T����0����a�=��<�t�)�33)��������u�����P�	 ��������c�* p�������)�\�8�\�����q���+����c���B��,������-����33�	d�����W	\	�r&]?	�fKKm��������>ܻ����kىٴ����� �'�Rځڴ���$�aۡ���)�r�K�~�����-;�x�1�y���.ܴ߳�+�]�����P���������F��&����ˎ��9�����ڌݒ<�����ѷ����}��b������>�T�V�_��������7�<�9�<�&���4�;����I���������� � � ��^����s�>���8��������(� 6�� lv_�F����Q�p�����|�$�����������t���}�E�������E�t���a�'�Q��`�e�������"�� 3��(p�{�ة;0�)*�*�+h,0-�-u.�.�.J.�,�*(%�!BJ.9�  �����o�~���������t�1����(g�f	�	"��׽�#���
���A���� ������������9���c�� � ����F�������������E��� �����H�(��a���%1 �"�%);,/�1�3�5R7�7�7�695I3�0�-"*�$�����{�&�$���R��^���	�h� ���e���33S��q�]��X���������YZI��n���������D]E"���I�r#�y�@�xJ!33q��	���.�y� ��`�y�
��������X����N���J�� ��h
52F+G'��x-��+�m
�>�^q`a�
33��pU���Oi�h ��l����}�\�X����.�����t����V��<�Pݷ�q܃ܝܿ����A�uݬ���$�eި���9�u���T�����-���Q��$���:����Y�o����������.�W��I�)�#���NŤ���o���ܗR�L���`��G� �~%
+s�N��t9�)�u��������������J	�����"�� ����	�������$�&p�������<� g�V�G�U�����q��"�`�'�)��"�������7����������D�� ����R�D�]����x�������2�N�33\ _ : �@������������������������������ 	       $ * 3 P E < 4 D S Q K I M S Z f t k ����c ?s^k�
AU_fjnprtvxy{|zxusqqrv{swz|unnoomjf]RV�a[bi33d�Rg�Dߏ�s�#�
�r����a�G�=�Q�������UG?F�	���7G#�*�'%�"�&2*E)f'�&�'H)�*�-E0�,�����y�K�R�    ��*  t��      Z�          �      `�      �2|          �      �:�    ��<�      ��$      `��      &	6	H	b	    t	�	�	      
d
�
          �
      "^��    �`      ��*          h      ��6      r�            $$+ . 7 D R ] O @ 1 !   ��������������������������  
  & , - , / 1 3 4 j f \ N > * + . 2 7 < B H N S Y Z Y Z Y S F ? @ U s q l h g  	       
   	    $$!@-@<@L@^@p@�@�@�@�@�@�@A/ALAgA~A�A�A�@k?}>�=�<;<�;�;�<d=�=p>�>H?�?�?-@  ����f�8�����������������B � � F  ��$$            ���������������������������������� & F b e M /     
����������������  $$      1 F ��v � ^�� -��� ��� � g��,��g )��)����E���     
��������
����������  $$   0 S r � � � � 6Vw����/!sb T�Q�_�������a�����.���3�����   	  ' A ? = : 7 3 0 , % !   ���B�����
 C \ I   ���������� $$  ����*����q���d���q����K� �������&�&�9�3��������� ����)����"  ��/���7�!���v�N�7�2�?�a�����'�����}���i�2�����k������j���$$    ����~�W�7�������������������U���X����U�d�����g ��;�7� S 1 $$  ��������\�X�W�V�W�Y�Z�[�Z�Y�Z�\�[�\�H�L�^�r�������������% � E� ; ��$$  ��� �x�x
�� I �����2�d������P�����9�w������ ���N���w�����U�  $$  ����P������<�����i�$�����W������c�,���`�?������:   ��~�V�'�P�v�_�  $$    - K p ~ � � � � � � � � � � � � X ����������   %   ��������   $$  ��^�Z��(�R�����7���������J��������2�� �.�����(���9���B� "  ��.��������Q�3�(�-�E�o�����3��~�K���c�����g�d��<	� $$  { g\RJHILS]	j
z����q�!
 ������]����6��h.c$ $$  ������B����������������/�O�w�c�J�8���3�I�T�X�X����� 6 � \� 7 ��$$  ��� �{��'�} ��%�j�������S�����$ ������_� ���D�����
�$�k�����    ������        ����������������    !!   5 p � � $b��0kkig<+;M_g`PNP�r   $$  � �tM8�v*�~� W P :  S����K�%�������Z '��b��� 	  [w�iXYYZYXYU	�
u� N�0�������������[  / n � � ,h������#�d�        T�G�,�Q���������������������������������

����\`
fsC	R�T�   ���������������������	6
	�����7���a�  p � ��6�P�� ��b utuuvvuvv�u   $$  ����(���K�F�A�;�5�0�*�$����"�@�X�G�2�&�������-[	�a�uM���$$  � j�*�����������������=F	�	I	��q� �&�%��l�y��           �vc	�a    �
��� U!#!K� �����o���    ����������    
�)�J	�	h��v; 

$�'|*�,�0b)�P  ��D�  6������^�(�����'�p�{�

����` 5� y|<��  
3���m���(�K�.���u��H�����=��հ�V�t�����{����{���  $$��k�����G ��HZ���S �"R%�(%-�-</�0?.�(�(
'�)G��+�i�_�����*�r���$$$�w� � � � * ���/����H����o���~���	'�
��
ViL����!�_������h�$$������q b