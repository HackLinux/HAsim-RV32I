Ǿ_DEսE�_�)�G����nxl�
2�]9=,b�"�Ғq�%����:�>F:˹诅�
��{��#S�����^��Gq�!�,��0������hZ�%v��>nTO�����eb�H�i���$jba� �H���F�}�|0a������]���`)�vh��P^'�o�Smǚ�qv톾�|�k�ㆉ)��-����'�@k�����f=/�^��<D�!�M8@�l.*�H��@0������o	O��}�8���fP֞�)�\K�m������	�N��f>(�� æjF����l�l�	<��8�t��|G���m��V��Q�T�=7u��F=��i"*��qH+�n *7�*�s7������E��v�EB���3DP|�T;̪LoWY�2�D�S�Tc"�F�+iq�
�=��ȥMU��;k�J;^���T���@�u�4���[>��ho	��v��+�΃.�I�쫃U��k�=��Ց\�k�/P��3�������L�q���l0C�k��#�������|>�bI�D�["ΰ.��Bފ3�v��5�%��%�Hɋ�I8�$m��#7]g-ܣ,ɓ�,70�u�:i��W�h�i�r<G:�y��c'i�ڌ�?}r]
�S�4�`���++;X����8���,S�M���Y����v#�y���t�����G�h�A�P4Z�u��U[{�}� ��-�l��r�}��,l�zN�sZ�F�X~+ɪ[�#�zm(A��-��n�Os:Zj#�j!� ��,>�̊���T1�1XÜ�zFA�q�K\��yً����N�����#طO8@'��f�v�c�jf�G%��Y��T�~���VG�y�r7]U�HUذN,U�8��J������Su�8BI96I�vkA�Q�a�[y{8ō��e�p�ҫ�Ȇ�o?��i�Qզ���%f�z͑�Z���>���}%���Ac,c�\`љ��H4"7g#�{��ZY�M��^��.q�m��׶�2C3�2�"뒺N��$w;�4��H�|��mSS�0^�N6qs�0hV.&V�.�ן�tk�S�1��~��˶�?E���? Y�A�"g�!��}��4(���l���^�5�Íݍ��H4�v$	����<q �|��1&s:��g&u���&�d�ੰn��5j��=��=�J&�_2hR���Pd��/J�Qd�(��EW�}�����4�bd�lE� A��n^ߖ�T�J��U�n�:��wm��u%~��TP�_�2?�g���Tj?Jz^&3���p��-���q�+!,�'o����؃����[Q^��*5�3D2btn���Ɂu�֒�>v$���Wr�ި1q	_{�y���e�>p��6c�ζȺ{��H�HƗ�ij7i��;�݆���ϑ�����3٫���k���-�dRd�iU���a�dͼp=.t��Ë�+.�3�;�3NPSPZ�������[+o�x���z�c�o+x]���OP�Q�SZ��g
�	�с�]Xpu�����ͅiM��CY�'�x��{��we����Y�"Z-��v�褌�p�[{�D&x��.X�x�:u��NL׾�EgS�&�p�Qg�I���F�6���"(m7Ù�x�ԯ�b|��\��5�|F2F��ݶ�ɜC�,-1W�������ϻq��d�~ە�Et�sr[���������eGeg���X�ηQp�������ٷ�v�nԛQ=&QG�:�4���R�`�	6��T�|����>�P.FO�r������5��:�����u��~`�(�uy��P�!�)3�8���l��W�P���A�nq�wE��{ʼ�~B�W����rz�a����W��V�*��b�l��đo/����颌��=g�%�"Q>�4\)h�OY�D�� }��*.�h�.��s�V�˒hSzxy(9���Qԟ������4�Gt&����_�u�0��Ew�,��kJ������`Yuߊ� �|���LtT��cM�0%�I2��0U��������d��a��SQ��뚰�3[Z��\X<B�!xDTO��B�B�э�i`�"@����[w�����D"���y$���6�77���&��]��D�`sIԿU�=<���QB3C[�٪�y��M!�g'bb���}�1�0���A��PR6��m��L�+�B�'���~4��f���I��'lg>�~#��bw"Ю_�Xe�2�"WK8I_�K-�εu#��ORM�,���vcp�.pe H??2��M��0Am���gԐ|�kk��&$��c�O� �F�Ѳ�rH>�L�(hY�+�����jY��և���t��UCmnz����ϑ`�7��3}{W��~˿��6��'��Ʃ;���[�Y���WaijՌD�m�5�,}4}�Ԟ�>�1L	�+��>U�A�Cx��o�k
��4��C���/K�����}���c���45��`���æ�:J��4F=���0U���<;p"b�4�c\ry�6}���z�f(\
��(����ha���/tG��[���6��~8����޶ 5�0���ٱ_�G4榮��0KD�m��Q{U��V�M�.����~Bz�O���\��4�Ig4~�ma��2n�� G��D��4�@,�o�J�$�:|A��������]��Q���E�p���|[�?n܅Z�N�T@��%L����A� bf]J�!U��m������s�x����b"��fߑ�?E��pI�/H:H���imQm0�h�q�lC}D�������Zb�������q.æ���6���z��A�c�w���c�M�%��1�����T�?����8��1,�.�;�5�}�%�dcdme'ߞ�Ğe�Z�X�w*��਒���}�`F��{��0�v:Z]U�=7�Ut/�P�4����G~/o	�|Sz3�K�L����ÚQ�.��ZܷZ-��)-=|��Na��/�^������O��k(g ��Ov�2W�d��iI7 {�lU>����@L���-ޣ!�1BF����/��y���J%Ɖ�g��?�������)�f�l�0�(��[���g��uh��߬�bD؛I@���w�%���%`R(倒Z���xI�oZ�6	�t�"�i*�Z{�w�/���_�"�2kbݎ�����*' y�n�#�	�	���J�����^=�IB�u6	D�r@7��E��Hd�#���������ڻn�|�0[PV�f�r���Ջ�|�[5��	ڃ�[o��5G���������{�%M�#!�p����$���CP�ϦzdS+F)[[��R�liG����<��]��4�V��7�'9Pf�+��ߏg�`�'�Jܸ�0R���ҏ������,![�"6+$����]J��U3BTkv��Rd=��������=)Ő
X���%���zr��t���\s�2������D:O`Z*�ᫀ�k����i�
b&�c�M@���S��{��k��lNJ �P�]��I�����eA�2�����o�)p;�5t\C�Uʤ~�`���:V��~�����ɂ?��J�Px�tV��P�0\]��H���J�=��d�n�9Fƕ��h�-��?�R�	[�>�ԟI�6�"=�3��ޙC�	���w��}e�Fu�s�ẹjU~v��B�e��7m�۷.�����u>���[���h�5N�\Q9!4��.�kE4�յ�ICs:�CEU��?�ĕ_��=��ԩD]x����J.$���}���ҍk�A�ъ&����}��Y���+���Π��d�V	�ɱ��-N�$f	/��8���p&TmL1���?MC�S5Xm�� �\Y#_�M�d��F��b0�(�����p�Q�\�K�C���I�y�
�d!���WFr���h��aޠ}�.E�f(��&����� VvE��s+0!�6���H�����-��g̴Χ ~	�kn~=�i�����q�[y���|^된4�42��jK����QBv��s�<ʿ-��<���P�E�x��γ]{��������$c[�|���g|�`�b�m�-�����A�Qɩ����ר����=>�Ћ�Bn(ҧս��!S�юZ�]�$y�)�F���c���3�-Y7���onՇtY��s��L[g��p4��MB<��)v1C�(^|Xdk��f��Fr�M��z�T�!T���;C��x'HF��^i�5�Ә��x�柞:"m�����b�-�L&�����Y�������3LŰ}���4"Yq6���gs��9��}��K����%;�+m��"cl�����x7m��!�_��;v�n��dBwCc`����@�63bd ~א-���B��5d��^&ŏsH�P�-X����"�j��3-$��R��+N��R�i{}�-�H�������_�c�^��Ƌs�U51�1�a � �mZ�ב�D�"��Y�\Y`X�7��ٌ(@�;�q�!l�n�}��*A���� �i����a:Ix�y��Iƞ��F	}M�sS�[�+)�g��k�s{��c��d]��� �qEs��g�3�,"*��y��5Q�{��s���"r���uK?��~��6��?�O��^��7����<�z���x�����|v]��{���m�[@R�V80(���0�U���NɑD�> �OK���@4!fp�E_�j�Rl�!Y~�f_YB��cd	=dc��v�� �u�ؿ�����(����|o�󪠐�\��uz��5����c�5�<�j���w��\�n���m��:�~&IZA\(O�������S!Z����2o5� ��Ƴou�s�څ5dr�!���	Ջc�/��9�BI9��U�BI��u\2.�k�{Bg�l�uF�IJ߸4in1�ѣ���y�D��^�	/u�$�Iq^�?����k��d:���W�����b���p�E~������;s�ȹ4�)G�!��c,{8D��+u�t���pU����M�(.�)"�9WT`��s/��%P��R�d!���)�M�2C F�6�I3��H>.���İ?->�E����7.��:Y4{� ��C�(=��|U��F'1�q���G5����-`9�yD�ˎu�BP������z���9纩�6u���K������ȗ�I��4��M�Ș��_�
�L�r���:�	�Pc�py��;�+5� �ɅCDK��"&���t�ޖH�بH���++�m�ߍ'a�8}r򘁚�+	%���d�_�Ԍ��uU((:��oH��qX�������ӥ�@m,�Wl�o�^Ԍ��H���d(��,��p�Ze��ʹ��e�\x0G��2��B@Y�=p�jQ�?���3���]�?�g�Cն�!����-����0�1.���TZ5��Z��=�J������(V��)D�R!��H���Y�:�Nzꮻ���fz�ї/L0ZkKR\́��U��J��"�C-��m����ݻ��&�xi�Ö�Sq�ܛ�J�0F)��2e*��m5i$A���M���I�������
�4����D|�*`h���n�xj,.5��R4%��F����߳�;�q�#Z��|	�4�����"��p�:�||ݷ�6�JK@]-���U�-$�!�N���a��T�n	���"��f��$Qܥ����+yﴝ �X�:���i�fi��!:I�
��h;���o����C��;+��¥���ׁ�𦘩k�{� �	�m�y������R���5�V�uC�7�ϛrn���Pr��ȁ?-� �O�>���F� �ƫ�0�w}Z)}�� � �n����**A�}a.�m��;�i�*j�*�J�Dw]sTT����!�?��[ʒ�59p"��E����}F�/I)@������IY�]���$��<�|��{8�������LF�GVQߔ�]JVc4�&��S�,�a��#̜J��b�����h{�Cʟ�c���`�Sm�曙�D� �:|uN�q��Nb�cG���m�����t�f�y���2��_ώ�k�>�?0T�9 �*�Q�r��_F�����u������2R�
��?GbHʖ�
����
l$��6E��O��|l�y�_|E�z���;�F��'?�)�Ԭb@���vd�1�)ޔ�����/�؆�Iq<�C{��w��7�nT�]y��tR7�Q�G.٥l	�!�w2����LÅ��k���5�Bz�U�y�15&#<f8����#��^����U��x(��2�#�]E�$�W�s��%�Z�Rzo)�z��Ҝ4��%J�]�k"��N(��R�)o6P2C7k0�GvFL�������<ӌ��p�طB��4�	o�TωS1�ހ]q	��A��Pb�ߖ}`=��E�p&�iov*�t�g��Jg���c��m"�b.�!�'�Lmgņ�ۆc.B�y��ݛB�ꮺ����X6�qS�+r��<��U�}ٹ����3�(�.�������
�A��W�T���FU?�N��1��~f3��#zP���[:^�2�=?�N�{�!Y���x���<��1�᩼�ہ�wd;z��d�KO��K�C�1�גx n����)�SA��z�N`$d�����$6�R���;E	e��t�"�<'i^89���n��	�N+��겇o�,'�\��'4�����(N��R�b��`:#��	��9����ٰ���4�o��J���ɐ����'�C��JB���dw����i���5���� ������
105�}��'+\V��;3X�1��_�{�>͐}���w:Zʡ$U��v�������}v�`�}+0R�N�Jb;�|�޲R��]b�_���d��Y�B�3{�l̚������
�d��N����5�#�4Me1�>�-î�5�/�գ,&dO�;�y��j��5J��q�c2^����1�3;������5�K;��}���D.��G��:���eѭ��Zׯ[�~W�Ѣ$���0DA=6<�ws�us?� 5����l��nD��_p�0f�є�j�4 ��ZݫC�XTr�^��D�z��^���y
$dI�_�#����5����`d���+RfcJ+������OLd�i�|�w6�5���yL���]ώ�;�n�����)f.~p*��g����FO6�X�=ɆVu��];9�(rF�� ��z�A�*�Ly(��-�GJ�{��Av��`cN�e^ i���g��C���g n�	��/�������. +�[���N�;���.wMm��?�{� ��O��BO�5�:I����bA��>jh�V�z)3n��]�]���=�"�h�ij�Ԧ��F ���Z`!u�er�.�?�x�SiDZ��I9���Cd��y���Ci���PШ#�[��lP�c��z�n5�aܠf��(S�BC���Q�5m)��-�Y6��Jm	��]#�Z]��r��(������	3�����A�dH�$Vl�R�͟q?@�UO��Q�7�4���.�2i�*�WY'�"q.ε�������ė~�3��2����5y$A�����@�a�Y�����^��-	��9�\�Ӌ|���%��%(���dW�hZ��Մ���0��8�=��ʙ-m�*>J�%`�=�dX��x��A,Obw���9�{�4q��l�zC��h.��kFg��X7a�G��Oq��eM���P�+Z�j��b�d�_ �i��m��qqb`��$�tG
n�����x����F����OMDN�U�}���A�ޮ���n�O���%�2 n�/X�1-�!�q�">'`�2iH��w�>ҩ���pr���i��i�a�W�k��{߬������
 �:��7Π~�\���[���y�������.�)")J��o��WF>YB��;��@9�k��v�➞,"?���z��d4��Q-u�(M�|َ�YT���S#�1*�\1�`�zL�h'�I����/��(���^�	Z���������Z_�僱����F)�9�ep&������P:����W�[S����Q�����zny�(=��X!�A�+�ecw�>�������?�.W2X\?#��5�>gA-ʰ�厣I������c$��S�<ϖ&�~�:Q^�~"XN�Fj2�r=&!�l-��;��&a���9��x������1|`i��BP����`rnZ�����e1�Tm�TB����1\��6k#(5ʔ[]k�T?	�dk���w?0�FA�xnz|:��l���`�Z�)�Z�YJZ�̋}� S��؀u$�!��3Ӫ���G�{-n��"�qH�l�<=h,6��m0��Ć�Y�jYωs\�گ���8��};�>	�+fΑǹ��,)��3W����t���<�6��٨�PQ�*#��i�y�%XӚ�b�V�>pC�`f���RV����>����ǴVd�F>ԍ	>��:pI�g�1c�W\�:%W1��l�R
�����O�<�8�����> O'��
"8�l>kp�E��D31���
����jt�|B���sf����� %]��q�%���Ҙ�R�rQLc��<���C�O.Y��yȘ���6g"0iP�O%����V��!ׯkBB`<�.]e�(G��t�C('������V���i��ǂ�b�����;�ٳ���3[���y^�郝(Y��Җ1��H�3��~l�Œ��ypY��i���+�3Ə�<�o&�0e�Ș��]a2^1(L	�)��g �\�x�b}� xd;�cՃc��kݾ$\V}=q��r[k�r����>�\�<� �޲�)
6p�F�)��<8�o����ݯ�
��s�n�,_��ëQ5t�/�� y���/ c�U-#b|h��!x���X���1EW8�XT�a)��A|!I��*����\h�t��&��O��`)�I)Q,6f@]őg�:5����3�͓S!,������0/1�\���*��=07Hoه����E5/ʛ��j�W'�fe�2��CruM'j�&�����hH_���<N��\��U9+YMA�Ҋ���`��~�u] ��p����*O��*a0͆-im҇
��U��!m
�[�}0��U��k��`�������=����GQ��="���D3z�I��Z���2R7? �v �]��ʰ>aF�o�&Ss�g#��[:���$�*�zI@���v'9��J"�Ğ	T�Zk��u��4�i�a�O`�0�����\X��$��6��u�顖��m`��(��G">#���o�6�="�lAf�1��	�!&�|C:L���;(Q�wU.�0��v�޳�]�Rҥe�E~���Z'�PE�!A�`C����z�_a��O�ٸ*oǳ !d<�8�m(D�Oۥ�@01��Jj>�6�Y��|U�f��A�gg��h�����K����'��"-E�����+�ҕ�@�o�/��D�v�EW�+ �� �Ï�04�V��@^�v�Kơ�NW�'�V[��tn�a����?&!����b�ޙ�t�/.�@0��d񀿾誼-���i���}+]��T���	v�I}MV�~2�k�"�M��p���j�%�g�v�Pڭ�^ҍ66�� @G�Ӌ6���4�e��lF�]"!����k�^Ѓ�f��+ʘ;�JzU/@�yv	W����9��j+W
0��^�P�tsWL�|�-�h��}�)S:>��q�^���J+cI�[��>�}�d�zd������}�5sh~f`��Zy��^���R;���]uY���T ��%� �S���������d��轤)a�������i�A��R��̮}�(1��p��"}�O󘭄��<��V@�A�"�d��{�eGvΝ��B�ǵ.�(�3�N�_]3@0 ���c�{�S2����5M?���|h�G�w}��tZձh��(�I2hG���둘�A�׹����q���}�R�����+̍�<��V}��i��C��b=�N�);�lя[��Ke�BT\D�ov�t���5.�����.��2�t[_R?&݂�P��JW�Ԋ�~e�W�46m�yVs`�H�.��ʔ���x�iF��e AB	�k����x�Xg|���H�����>�����O�'^hL����K�0�����\���-mmȒe�zBc��Vj>�J�tW$^�aـ��P�����w��}��eMDu���`�h_�����K	������pvl^P0��"�0@��ٷ�� ��`68�����C�to��ʂ�gg�㯺�)��0����<E��Wg���ކU�%Ws�E��
�k�k��ڛĊ��.�	�R����y�\o���ؗ;�.�V��U�_E����퉋� R�IW�����y������K��:��{@_c2��JQ���푱�C����2�k-
1�qP"	���G��J ���m�S �L@��V(7���7n�i�J��6�T�h�w7�~R�19�~㩧?�Z2e�7��t�]u�-�P�ჱ�J�(�=������Y'#������TG>rLи�է�*iS��ɴq��(���x��;�P�@Ͱ�_00_���ϒ�h��#㱤]�,��/:��/��I�~�x8S�|�&�H�����eUbγ���>�H�G �V|t ���J�s�|)�%�2w�'���j���Ye���綛NW(K��pa�]�]��I����w�@��c�l��#��d��ym�=��E�q��]��\�e��� �x����(��$�}�J�a���m�1�{�=.@�A,�}�Pse�l7Sk��L{�{�ΤN0!�!��t�����H;��8��"�dZ@}up���R�M�����,Z�O���.g��1��v�	*_���ѩ'�d�6�f�uhZ8�G���M&P���}c�\.�� �i��� �骦ј+����	��_�ӏV�k�~`[|�
�4^f�+r�?�	���G&�D����t��9x<A���Ȭ���&|){;Õ����x�_Ϟq��	�Ve�Wn�V�P����h�N�vI� ����� ط�RJ�Υ�#D˦�T� ���#R�k�$g�i�Nҹ�iș%%6�\��KR�����<�u���&����ɖ�;�WK�(WBO������vԩ���� y��g���>���u���4Ξuʿ��P��̀�-2��-g���X�������U]��,ςQ��tLeC��1��u�>��µ���$�.p�(�e��(3�gr֯t���᥋ܷ_nnn��<�Z�[�A�V�� T����"�*�)Q�w�|y��V�հ��$l�K\���ul/��:\0��kyi�QS~T�:�!�`��>_J9!r�hT�i���I�&������S�	�3�V�xar8z�2[^�v%4d�wr	E��q��bS�5����	G���Z/�+]��[H�깊T#�'�G ������|I&xnx�	�5��������\Im�����a����M +P$ީ2��L��I�Q���:�s��瞸>�"��0��`��] �InY�|,ɣ����n��or�m"�%R l)����:T�)�<\l�l�O�Q#�����S�" ���w��Ͻ,���ԫ,��	Eks�%��H����<1Z�	"`�I8(&v,�>�S������N�� ���l(�HԘ&��S$`v
�2Α�g�O���o�	��k����Mf'3C�N��b��bKO���6�s��(���!e��ѥ)��.�;t3��,\j'w%غ��-Ė�MJ(&Kx6�R�>��Pϭr������\L/�#�M�kJ�!����;��]h�#�;�	���LSj�0{!B�RGh��kU�^g`O��V:�"��-�~�Z@�*���//��`�K�Y!�(DH�4�{^���U��jxQ�E#!����a�_��+8g��:����"�ȹ�Ҫ�76���rP�_���X��m����E���r�[���Ѡ�<�3�c5%�=(%�GAHl9_MOz�J��o*q��R{+������F�!���5nNK�3`��mt�0����2�RԴ:���9�]mF�����j�ER�u#�?��h��I�9��c��y���N'>�tB$�����ZÏ����n��c�瘐\40��Z��QB9�+`��|��H� b3{>B[��S����̼t4u5��EʕaE����:Iǽrc��}z�Lj�݌��MU�i)��(o�;G��8��C�*E�p����>�'c�Y6`�g�#~�Q8�
A��?�T�)�f$)�=-�w�މ���.��O�
[����H���p��+�q�Kl/sv�e۽��?��Y
9f$M�WCK����vD7U��R�Y�c:''j��R�{��	E�*b����N�����h����!�� A
2�6��k�89ҍ�����3�H�������ͧ�f��=����Ýt�'tOťZ�+b���yV�2(����}�.]ylHB��*U�h��\��(�_��5)���䫇@���7l�|>�tN�C���y�����݊>@��{���];����.NW�.�,��vEy6�67C�������>`۲'�pe�u�����r)�W����ފqO#-sp�}�@��4�09��A��cc��ζGtD]���E����G�F�1#�}ظ�=J�@_�vc�p�8\�$��H�O�T]ti�
hQ�Q��a�@��E�q�4n���xߔ�3I�!�d۸-6�n������q�]OqL��,?;�L^1%���X]�ں��$���A��:фٌG���}��!E�얅�uo�]�zG�3��gx�*#B+��y�e;�W��-	�!{Ϲb5��vj���6�8��C�3���Vxm���S�@tW	��'yd�x�k���d�r�9��T���� ����VSڃ��y��й-j߳k:��΋G0��<LF�Eы�a�WH�V�H_�᰾���?Q�.��m �z���Q����ӱ`)[X��93��s� ��4�ʓ��L���:M�
�ø��\I(�M~�޾b��-�&�cm��rd!��[�:#�v6����'��M1*X>7�J�#:cR���pBN՝�a�5%��h�L��u��S���9�� 0��؈��J�
�+'�������qc����-���F�:�]����9��TQ"�z]���T�����~>b{Ja��4mr�TR.'�2c*16^(�߾B���vXE-s"�4��V���1t��;��\���r.FቝE�_|���鍄��?N�I��貛�F��{���]��iU�L��6��7��	J3h�>�����%f��=b�lE�[Q͊��҂cJ�O�F㪺�"�*�%a����S���\����ï�vupzwWw�xg�7���j}y�1C��l�'*�)q�5A9�00�	�쓔r!
���3�|4@��,bB�?ޫ:�o������'��9��L�����Ɂ�����c��e�Z�ˬ�{I��p�}����*���V�%�I%2���Q\x�����Y�B�N/�@�1k�g��1E��./&L+���CU狕��k��Y';e���	}WZ�
{��N�m���B�uW�%�p#�[��̽r"��/s�
.�w�2��I3���d�������[)�I߼f[,�w
��%������1@d�.i�dS�em
���u��"����Ş*���z�7�=���2jr�ν)Qd�g���ˠ�wZZ�[��4�ᮄ�`���
�KC���K�;%�\I%e8�b�,�����X����IU�` Gن�?�����d�<]��F��{�}�[�$Z�3���D��G�d�����y*Q��;��h�$#��i:�~Ќ[x�օ�ႈ�X����4r�揌44���X��x7w��#~��p$���M�7\��
NCץ���#�"i�=}7��@gu��c^{$ƱL��>ݕ�����FE3ޔ����}'�\!��1G���	(�`5��hKo)��U���I	q뀥�F��l��/�����fU�Q~�_�	E���p�0��*��v�K�A��Q�)>�hJ��q�� �f"�S�гI����H���mh���N�v�I�t3F��ƙ�õ�4��E�D~��s���}������k���4�~���l��sY�ra���s������Q��?���&_H�e��<�@Sc�:b��z3��͐-d&)Z��yĸ0��[��Rg.n��b�,&��ϋ�Z`��`����<������2�$W�S_&�+��2�#g�hl�Q�P׉6�쥚y.`���"��I�����4&��Y����^�~�aB��M?ob�MxC;^���X�m(1nD<���sZ5�H8��QmY��RC���_R�]��N+���Vn��vm�3�H����C� ?����fnE�dcOo,��5�(X-��o4%F���.��]�W=Z��Q9G�	T'! ��e�����h������c�������������5+�-�=O�=�UZ3�͇{�ݟKZ|(}¡�#U�:q����f�h��������<F���DZ����P��s�����;)=)�έ��G�YJ#����,ߣ���I�����dc�Jd���L(g�^d��^��I�q*yS`ު��v� `���eC �|��ݟ�M�Wt��l���m��J�p9������0�#����ĩ�ju�a��4��� cz��qC�qc}��cũ���f��9�ؖ��� ��bC^����X�3pn�mfUD�����i	����gH:��~k1��p�pc�������H��)քn�%����;���d����b�������-����c��g1좧���oz<�������u��Kj,�B��}��5 
�;/cn��_�E��袑#����+g����Ճ����Fg����c���h��:�l����������M&��T�c����兑
����B4=���&�Bp+0��5S+�,*{�.�vB�X��پg���
�v�w��Ը���suwdf�$� ����p-���r5���Xԋ;�8_'��x,�^�(HddQu�ц3�VE����Y��0�$�d��q�:�}V�v��h�Y�g����D+���PK�g��ڃ��y�v�$���踤m���(?Q�!�0 �������U:��)8�b-ؓ���ӄ� �҅D�r$���aI�c!P�C����|�MV��֋{�(ȟ�zmd�<l��������,��1u��������!�akA������Ɉ�)��v��DC�(Mo��+J�����tL	k��-5޲>�[8Mz��0{���]�6�L���I�x��犓ujy���L��C�����,|f�k�vg��G��l�daŶ����˨ꡡ���r�
�����*�a�@-��5�� �����rA.������6F��6>�$>��Dyô�a�/�wi��ik�j N�P���k@�c�Y����6��V��!�I�(���Z>������=L`����߫�p՞��~Zތ1ݞ8.���,�'�<�j�Y��/2��Cj@���C���y\3�U��h�{A����L��_٥��+6L(
�������?TQ7p���4��I�+U�2>�J��b:������i�t�z.jF��'(��s�-���@A�4
ث�~�ʞ&�+�9��^�s��Zn���z�M��M�8�՟�V$I��c �������s(�����P��M|s��5g����(Ї��E�����Ol�#>��+B�4j᳠��%	c�����H�E��eqH��I���5�������2A�"-�C:$���򟊝^�`f��I��9�B��ٷE��bR����%�!�6F9�	�D7�����0P�����cs�2�m�8�b`�,��ͪ\3#�9�_�@n|	�,.>��7+���uXj �Å��^�n޶��@�@0F-ִ;A��dJ��в1�6B�q�TN�p!��r��ג�C�)C�������cO3t�ew{�����8��N�rA�3"
��I ��o��s(��a~�h�����b��=��7?٬/�D���� ��W߼k�Hb�|�U�\������������,�A������)�C�L�)�xOኗ��z/'�<C�޿CR��`?`��!��m���ۦ��@J:t�|����(}��}S,DC���JQ�M!���(��C]�a$-B��r��/�_������Bm\��>�����m������>K�4�gb��A�0�bX��!p��ue�����mq�KHQ!@�/���b�h�9Q�u�%k����M�����h!ڴ"�EK��=��&���{F+��Xp�o=|\7ޗ5�0�/��8���|�����-o��\��P#؟<+Cs�Jxϼ��L8�c������fl��M%���/��7�bl���P�u>C�H��A�r�<�����	f�eg2��Z�����U ���Bk:������X����e{�D��vf ")���y��-���f����_�,Yqe��0q�Ѽ��Z�c$9��F�e�;��f5P� ����E�ͱfo�'����5N�:	��r $*����|����b�ad~�KG��I��i����U��FA��|�Y��e�S���#����g=Pj!D��=Y�h�7�m��<��c�6v�l�k~mæ��j֓Fb�}�r���噠)G)��t����K��~������֨�!��K�k_G�+\d�lV�H����!!p0�?�(�w����M���٦u�[�n�LU�h�v��o����V}�2!+��u�5A�E��}��{�K�FRq����{������A3�U�����䔔R��8���+����b ���Ad��d��Bڬ��X�g�I�k؅����y��(�*MrK���YR׽=9�%����5���*�"���}�M�"�%s���/n7+�A���Zݥ�Arh�ڃD��;� T�m�%������?��^����8晩�E�/%�1}���=�O��,1ВPJ�gi����䓠-���r�j�0�4�v	��]��]�F�0Tz*��nX�8X]�	y ������5�B��U����<�>���#mjk-a���c�)�PjWnkhmniHo.e�H�$�t%(���r@1����6{�l������a��|��׉r~׊Q�	D#?��Gꄤ2e馜@���gU-��2�W���9��3;"3^�S%��z�l98�?Ym�3���_QW��e�}���J�"���M���[]�$4Vcvϡk��0��y�}��T蕎�����G����<�<�֡�^Y� M�(�Z����L`m�3Ǩ�T|�(�����ip�|N��0�p����a��ɉ�O�J�)�Q�f�!�k���lb'�:�nʔuV�l6�>h<w������yQ
�쟣�ݭ�{H�|4@�e%'n�bh�tԩ��4�>�>���k��h�Qu�4,������2n⥶�_�����NU�\����
����^�ܛ㭦�I�梥#kz�rf�j�z����*���-�r�gT<��e�e�rI�b`|A1*��
!vӧ�"��K��^�������c�Z �
����{�Q���	틇
9�[�J��K���R5�([f!u�	.�����CF���m,�J�UAw�e� @^��1e�;�m�v^�Sf�ǯ��l�y3�H���ɞ�$Nk���~�>y�&�T |]g��/u�vD0��\I�`X�ޓ�� ��W����_�$��j9!�x�BCf�w����󞭿���X&�z�ࡎ��W���=�cQη�E1�md�ǳ�o�bq�Y��^c�h��1Ƣ׾�\�����^+��g6N���nۣ{{������g�.!��&l�Kڔ�&+�n�~�i0ǫ��w_��P�&��`�	��� �v�3~�"7�Ұ��D'��L������� }�c��.T;�X=�b�B�M��ݰn�HaU����z���d��SK��t�wy�.�8<��yǎ��Wٹ��AtMߴ#��<��Y�4�;���0R����M~Jr������S�!�F�r�(�U(�Ƴ'�U�n�� ي��v��`u�;⾔��%�Qw����=��cXuP�g�V�}s�E��T�����e�.T��S5��k�T���|��݈v���ݱhSL>q��e��E�ᙾQ����Y��������4̙h�,m��.�.�8�;|��<�u�C��vC�,f�>�V.�:i�f8�ʷJ�{�k�L����U
�=�����}��a�t����o�gS]M�88�Q� �	�!R|Mћ�ܪ>����0d�_�˥�-��yC;ζ���������$�T��-p�2��D��jb����ϣ������������U������(�(��.�[c�ͥ��G;U��˺fë�L�&�2��L��� ��$��4��G���Ƅ��i���C��L���b�'i�m&��L����)�u��b.�r�쥼��v�f�lŭ��v3;Bf�������7dG�a�����6D������)$�HDͼE�KwR�"����Ep��!VD��������/Klyв�6|:^�b�gI�#3n�{�.����B�fC����UZ�8HC���1m�3�&��ʴ�QOe��fz[3���./�Z[�Ѻ���>�'#�����u$3��rAL=�J����ɗ����+\���?fZwt����'jԮ�*&Sga�9:"w�
|�
�j��u���6LŦ��]�E���ݴ.[($����pD�%_3c`:��7h�l|��-"M�VY����\�C���s�	#�%�e9	S�K�:=�?�����`zAr�%�:��@��j�-o�%Ly�Z`	���y*\ɛ�k�ozy6s��#*~�,�p(�_Qݠ}7W5��+���O�zL�$�%�������JA����k��.�b� ��>*w@�U�-��eӉD���yŽ�h��2���'��$�E-�����˘�&ŀI<�V�c�㿏��	�ӌ�/Pu���o}�x��$�fc��k�^���J�
��_�Y|xS��߮�ABH��4�M%X�>�Y��5C@�H�0�)��z���T�~ꃿ,.py���W������ARo11��3\��P��m��٦(�R��-��Ć	�^���5��wv+G��h����C�8����b�{��}Ң�)1��|�"zǆ�gX����5Ƴ�{y�l#Hu��e�"�u�`N�.�+�t^��(E9ö�p1g�Fx��im�@�;�Ӥ~37��ԁZ�|�#��.��7=ߵ��o2U��|ٝ�^)�*�RT(d���:�+�0��IL2��ܔ����O�O#���^+r]LA��w���=2�x�͡��pFMF��lW��(%3��5��h�,��b:y+FS��&=Q>UR7�I�U1��R0���Js�=p���"8�:̋�*}a��9[������i��8DS����;��G��oe���:T1���\���5�{��t/�N�u�ra�9�U�wq�t�F}f�Q(��㤕�b�VkJ@�oK����m$�w�G�8��GR�����c��O2IBB�Wl`�_ ���Ǝ��0YFUk���!�
t�0n��19d�b������38�2�u��Hym���i�|���W���z+9/bޖ=���s��6�{��mR.Y�k��ҥ6��N[�69��.
P/E;3�Dِu�dG��4�ʀ|�=i�Cz��jޝ�ʜ����
	p�*Ȱ���~��YA p�4E_gM;o	���T�I:����RU�f�����X�U(�d�QƄC�p4�>��5�)\;k�A�%���s?C������* M����Q�Y��l�B�f��i�6��;JE�)j0YI �T4^�D^<�������l����b���&����e�Y劳�e��}3��fV^��#����e�Rz��,���H(W%��>i��s${ԁ���n�3�/������7'9?ݧF�e�X��:��g���9\�L�p\�F�-�������\���?�t���jy뜊ӓ���:>ŧP��73�S��3��Y�����Nc-=��0�䔉'@��ޘ?;��	E9�e�8Uk+��I���)�����s��hm
Sч;E����b��F֏�pCѫ�,���}�,ŗ���K�	=�X�ツ������j@Oo;g)*��;r��(�AҠ�S�}�k�{��� �Z�vˊ��o�