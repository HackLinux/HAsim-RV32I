��(5ss����Ԁ�U��h��UB�ܫ�� �ݠT
�UHZ��M 8���­O��8��� ��}t
���Gs@+piV�o�h y	� SJ��}Ƶ�B[����@
�
Y�O!�o�	RC�$ۦ�I��>�����_�@)�jX�s�7�	=jG�q��u��Õy��U��΃T
� @�R�S�{�$5�9� M�Qʟ%A��:�� ����@%A���Q�����QEEhG×��}?�V�M �?ܯ���@�ʪ���zS@r�hTF=Λ�j�up��>b��*��
���3Z��4 O��J�j������
�U�Bo�8�'�G�8����5�i�<������(�����:jaOJQ$8���:�@X0n#��7��2ԫ�j;����� ������!9��5p ��*��p"��DT<y�h���8q��EaʤFzz����>�aۭt ���?>?�j5 �~�/�*�mAMP ������}��!5�v�n
֚�����(�BG_} �o@TI�s��j�;q4
�W}������EO�n�	5@
jK��@	�#�Cǟ!���8��U
k�;�TP���!U��5@�P Xn��]@+�Z�%V����CӅ@j���@p	C@���5QO�2Z��F��6��&=�Z� ����r���ꃏn���	;�L ?. 2�?����� ��d)U>��R�����+QĠaE*A�� 9q�)��;o�r�׋H�zсDW��2Ui�gaM�AƝ>5�U�� �*(�8�xu����o��	<���<�P
��<xs��������r�� �:�8s���6� 4F���Y�W@+~�������� �ڄ����Һ 
��!�q���4�$�c���  j\�>_�uP��ƴC�Tv������$S@$�0RW�q��zj �MT�?�b#?~�4]�h�_�;�|*	
A-�p5�;n���-N� �W���-Rc�h���?�:�$���|�^<�Jk�:� ��e5�㾀4#�F)U�s� P�W��51���	<���q�ܒ�����*W� }=�|���p]�W}�!�Q�v4Z��hn��6���m��G�x��O.cۦ�Ó��
(��W}@,r���P5�	�?�7%�����x��r�\Ƕ����S��7�@9��ȇ 09mP ��A��O����Ù���m�����P�P�]�Gr�q����j9չUy�� 
G�re<j�ƀ4=@�{���."\�C�U� Q�w���Z���Cr�/NC��z��@$ra��U~'��o�K��C�߇���	�ۛUw<�m������a�c��F A��"�K�)�@w]�`*c}µ��q��7�
�ʒ5yPrj�,��!�@QE<��>j��aˋ��(����F�^-^F��t��N�H�%����k���1�w�i@p���2�O�5�@p.���o����v�<[��s��u]�hǩp*����X�D8a���n4U��u`߼�h
߇�T��r� ��S�9�� b���@w�� ܾU�� �ҋ���m] hO��|���\d�)?j��
��@��}�@R����U;��@)Z�9-@BMi�;�Mʚ�S�v�@T<{�Z'�T S�8����t�n3��F��`!iF�
8�.��R2Ɲ��cS���:�P��ӈZ׮� ��NM�Pצ� (P�"��
���'�o��%�om ��_�o�ʀﾠ�÷��Mz{i��-�%~R6���Vܷ��7��� ��4
@S���������ہ�i� �U�l����u ��BW�U߉�5@ |xT�*w���ǅTT� H
?	O�A���۶e�ǥ4/��l)Qˮ��`�k�b0�^�բ ">"��x�:��S I����1��H髬���( Q��}�[�BI��'�CzL h����^��h�0<(Cq؟]0ڼO�Ƈ�S@u��hw���~5���� 9q����:�A@{u