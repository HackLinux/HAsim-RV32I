��VsZ�������� �Vfi��5�a��9R",�:T�'^�N��AsI@��8c]�l���d�Z��ZZ�����xV(�ZƋ�[�6�4Z�##�B�}v���m,8��^�b�A+��Z��dg;�b���θ��܇��`_�'ǥet' ry���b�D��e`]�\zt�2�7�b+��T�K4?�X�'��=����:&���$߇�N�]diY'�$���J��q��h����w��K�ȧ3}��E�n]��D�Â7~���-�8���p� ^�r�,/% I��"��+��wv��'�_�~5������t�چ8�'�G�0����a򞽆��hu�/W-�ոG�|6@4�S	�~�s+�Rsl.@�ɀM,��C<u�ι:�Upv�~m!߲r�Hny�Ԙf��kj�v2����-3��P�_�9��!��9��L_��Z����?�(���Lt�#������|���e�v5d��6�-��2�L���]�X���,h�T�e�Qc������E8��;�0��&c�=,�ů��X悧�y�2�!�b���#��D��bS��J�Aj�'o����/feoȣ8'��+M��"������G�r ]�5�ʾB���拹�f��A���F�5�����o�U��9�&��8e>�¢��м�KS�b��q�"�����_Z��šbb��)�3VaZ���ĸܣ�V�D~|�1�����3�
v����i����iy�U\gk��Xeo��k�&�C

C�o>�sƠ'�2�VB���ǅ�#{�x[���e:A���#�UE�~εql'S	��T�Z�͉�⁴���vԕ�]���|KƲ$�":P�1��6�y~�6��^m4J4��8�#3�
�W�<F�߀ѕ�3i����x���ӎd{�0�e�U�Dz8�4͊���#�v*u�j��.su��������I��-�B����Y�������������OD�.u��$~�QMѵ�[�'����3tWL>O�.���c�z'z-������v�`�1씶^&�>�k���V�q�� t]P_k��\]ן�.�]ж�4}9���s�ļU�����"2Gu�O �.<aō��CG?���Clc{��wI�,Ԣ�������B�V	������ԝU���-餫��z��� D]��.��*ʃ�ᶻV "�(����dj����a�Vpa������Jo��o���iD<>����e��$�oJ��7Yd�Q4�R��Gpu��cr�����z�f�@*�5�H��o���1���i�����W��Vd����j�#F	ƚ�X�9���F&z��9ɪ�@�č�V���`L��^�U"�4�%
S�&�	�kl5�U�h,��v�w���dy[%oK[���RHy�x��W���jc�\C�F������7�}��!���z��x+� �Ε�%��d���hh&�o!�m��f�A�-�u��H��tJt}�z5�В���[052�q��Q��Q�`<�+�EQ��x��;��F�k����͔��E/vNr���>�����܀.^��Y�Uk�@��)�����/�un��i���ae��2��ctl�F�:qOՎǓ�@*��@��eY� ���¥WlEn�~ص#�Y���w:ţ�C����U#��'���b\�dTd����G���o��%�4�/{T��۫���@9���Hm`��7�u鬍���3W��&c�7�/ȕy��|���#��A���MÔ�����]<�=Ra���df�5w��D�:�S<�����ID����ǉp׾RP�k��y������v�m�;�ȃ