�������������������k���w\����u���������-���������ѽ��������潈m�����a�������������������������-m����m���fzhFMf�������Ld��ܗz?��槯�dDGm�����k@����������������������������������������������������������ad%\�ĝii��ug������>{�������������������򽜂����pa��������������������������)?f!'�������f->>--C`�������s���ƃVDN���@$.6$%@+8�������Ս����������������������������������������������~����@w�ʝk|u�����u������`Yrz���⽽��������������_i������������������������������~�pM�������́`FM��Vfm����ѧL��̰��m,L��@$n�k��������������������������������������������������������d����ĳ�ã~~m����ѧ������z������⧢��������ձ���潋I^__m���������������������������u�ud<m�������̗z7f���f
2M`f��gd�̰���]+6����k���������������������������՝����������������������������W������È�uu������ࢽ����̰���������m��������������ËiII_mp��������������������������~WU����������ƨb`��܁FF`����um�������OD���������������������s�����������������������������������������N�����ϟ����y����⟟����̺��������ua��������������Ëli^_V��������������������������ʄEn��������̰��{b`�f
m��Ɨ��]�������ل,������������������Ѹ�拯��ل��������������������������������������W�����Ѱ�y������ϩ�����������������gN��������������⽋ilIAj����������������ǽ��������۶�~�������z����F>-
`��̗���uu���������m������ѽ�������������|����k�������������������������������������ʝ8Q����`j������u5�����������������g~�������������ý໋_^0Am��������������������������߶������ܗ����z>11M�ܰ�����V������������������������������I_�նU��������������������������������������}/���fV������dD���������������������������������ýկs00)Aj�����ѧ�������������������������ƃz��ϵ�mFz�`!5M������Ѹ������������������������������_d�ʳd������������~��������������������������ߞQ8�������������������������������������������򝧍yR9))A_���a���Ѣ���������Ѣ������������`���廍m��їf5`������������������������������������௔ʯ�U����������������������������������������߳w\d������d|�������������������������������������uyuV9&00:3D�����կ��屢��κ�����������ӗ����ԫ����̰��PM����������������������������������ʽ��ՔkWd���������������������������������������߶���d����]@�������������������������������������󽧍�f<900:I]��u��k���ǩ����ш6���������Ѹ��ԫ��������H-!'Dd���������������m�����������Ѷʽ����kd�u�����������������������������������������}�������u,i����������������������������������������u��ffVD_~~]m��$6$:����̰��̽a3���������ѻ�ʿý�c<)!-`��������������������m����������౯������~��~�������������������������������������������������L��������������������������渗�������������ç��f`c]kkdVVa,$a�yp��̰V?GG,�������ý��d_�ԔjjR9<[f��������\�����������֗�����������чk���Ք@�~L�������ѽ�������襶�����������������������������~�������������������������ע���hPhppp�X?V?���ѧmF?3%+Ud]<3G~�����f555I������Ld�~I%dL)R<9M�����⽽�Զ����������ް̰�����������~�����~:@�������ܧ�����k��������������������ѽ����Ԕ���������������������ީ�⬢���tXPB(7BX����ϧmD3:U\U3)_u������F-`M<)�����կ��Ä:D]RVf������������k��������f������������Մk����k@&LVVm���������␽�ی@��������������Ѻ����̽�����u��~�~]uud]|�����������������������������yXp������Ք]6d:]�������m!fmm���f��ѻmD~�ʶ�U&,]�������������k�������p���m���������}����k%u���������������ʞ@Ud�����������������Ѹ�����۝~]D$s�ï�~~�����������Ӻ����������̢��h�����w\��UAD3&,]�������<!m�������zFf���j)]sd��\ 3�������������������◟�Mm���������}�����k%8%]����������������k8+:d��������󽟸�������ޟ����Ꝅ��d~������Õ����������������������ΰ�hPP7Vdk8/8U�����U,s�����s2m���ϣ���Ɨ�����]2auU��3L������������ձ�����Ӹ�z������������}����dE@:d�����������������:&+Uk�����⟈������������������������������~���������Ѻ����������Ѱ�z����~����ĝ]��Ѹ�a<!Ks���_2m�����ϻ�°��������m5����U'uuL������������⧍����ް����������������ϧ]k+\u�ޗ��������������L%+:~��pm������������������������������������������������������Ѱ��̺���է�����Ê����ɗ�`!!!������������������CxfVL3D<?�ѯL������������̧]~�����������������ki���udk~�Ѣf`������������UU@@%+U�ψ������������m]�������������������������������溩������̟�5����������������������̟M5c�����������Ѹ���������Ɂ�M5]m�����杄��������̽����������������������w:u���d+k�g�ƨf���������~���iUU::@:%D�����������X,�����������������������������̊���Ӑ��pm�z�ָ���m�������������������������������յ��������u����������̸��d~���������������È��������������+k����L@Udy�ƚ�������������i;L�k%���ѽ�����m5.a������y�����������温��ѩ������������Ɖ�zh``ff`���������������������������������������է�����������ѩ�d~�����������������␽������������ø��W+:U@%D̰�h�����⽽������kdgu�@��������m	!--!V����������������������������`rz������h�������џ�������������������Ͻ����������������������ѽ��]����թ�������������̸��������8�����kW�\����f��̽��̽�������ญ�\@�����u.*PH!!MVmm]�����������������������������������Xhm����彭������������������ϸ�����������������������潟��������u��������������������i+U��ïng�=++.���������⽻���������öO+U~��?mya*"7FXVV�usL3_�����������u�������������������uaaV?�����Ͻ�����ѽ����������ཟ���������������������������ѽ�]������������������dkU%@����gg$$$$��������������������ѽնk,V�������yG<**MPfc������kU_NLu����橈���������̸����󟁟��V]VG?<V��ԫ�ϸ����������������Ǹ������������������������������̟�ëk�����������<'',\��nu���4#6*u����������������������ϔ�~��ܸ����Ӹ�m.!*Mfcu������ddLLDLDn�~��������⸊������潟������a?4G�ի��ѵ���Ѹ�������������я�ɽ��������������������������,���������ѽ��a]g~~:%\�����ћSS6#]�����ϊ��������������m������ư�Ƹ���P*"7X��jsuuumug~���d]~��������ש�������������5p������a#N�ϫ��ϵ����z5,�ɧ�������ff�ɽ�������������������������m<u�~D_�����⽧������ÍN'3����ǩ����e6~�����.p���������������ɟ��̺�ư��zhf?*<f���cm�������ѽ��������ѽѽ������ϩ�����X�����⽐S4.�������ϵ���MLNAd������������Ѹ���������������������ܸ��ո�p����������������⽐m<#L���ï�����W3���$]���ɽ��������൸�Ѹ�Ѻ����zfP7*,Vp���������������������Ѹ�����ս������ї������y��eNe�������ʍXM.6$L~dL~�����������������������������������̰�M5������������������yGaeu�������\E=$UdLddl�����������sm���܊������⺸�������������������������������Ǡ������������������␐��e�������D
LLn��L%+U�������������������������柁�����̰����h������������������ѩ���y�����WWnv�~WU36d��si�}|��LLD,V�¸����p?������������������������ӽ�������������ՠ����������㢰�������⩴��������U%=~uy�ǻgL@8�����uj���������������Ͻ�����������ї�f��������������������̩�����Se���Ð.6a]]s)u������ޭMMV��]m���Ѹ����������⩩���������������ཽ���۶������������������������۾��}U,Nd~�������⧘k&*V*
����������������ѽ�����������������������������������������ǩ�Xy�̊mmV99]����h������������������������ѩ��������������������ǩ�����՝k�������̏����������͹��\Gu�������������ۄ$?*
'����������������Ѹ�������������������̰�������������������������ѢV�⺰���f����̸�����������������������������������ѣ�������������������U������鰏������⽱��à�W6]�����������������n+NaXV5-<���������������џ������џ������������Ѱ���鸗���pm�fhf��������������Ѻ�⸟�����������������������������������������������������ս����������k~nL��њz�������є�����~u�������������������$=N�p`�M]��������������̗����Ɨ������������潈����̺�Ѱ����zM?�������������������ܢ��������������������������������������������������������������ꔀ~%0R�z��������Ôamy~dg����������ս�������gg==�y���V<��������������Ѹ���������������������їh����������ư�������������ɽ������ް������������������������������������������������������������WkiOO<Kh�������ۻuGA::d~���������ѽ�����������vN��Ѹ���������������џÍu<7`z���������������̏���������������������ϻ�����l9���ⰰ����������������������������������������������������Ǹ�������ѩ.k��}_�����������կ����u�����������������������v��ѽ����������������dD3,<fbYH`z������������渨������fM25mzzxm���˻�������˕s9Kfffmm���������������������������Ѻ����������������������ް��������m~�����à�v\��������������������������������~����ß����������̟����LD]���Y`zz`M������������⁚�������ɻ�������˿�����ҿ�ˋjjm���s]VV<a�������������թ��������������ս��������������Ӹ��~~����pG�ʫ����k+Ev��������Ѹ������������������̢�~����~m����������ว��d����޸���޸M7������������M7���������ɵ��������ҿ���ҿ����˻������uVa�����������]aaJBTZp��uu����ʠ���������������̺���������X�����ï���v���������Ѹ�����������彽���������k6�������������=������������ш������������ff�����������������������������ҿ�OO/w|~,6$$$::=k����L3$#4GJSn\W\UW����ʹ������������������������y]d���՘��������������ѽ����󽟽���ç������������$�������������3���������������ށ��������柗f�����������������Ի�����www����ĖQww�Ğ:E\kWLL6DdudLLg���\+@\v������ж����������yZPp������ѸǀD���ՍM?y�;vv������۽������̸������������������U������������_���������������������������`5M��������������������ҳ����}���w/w�Ү8k��������usau������v\8\�nn������nup���pZa�hXDus��y��3�ϜV*7X���ݥ=q������ï�������������������ɻ����U~�����������:��������������������⸸�����cf��я�m������џ���������Ŀ�|��������OwQ/\����ʫ�������sd���ʶ�k}@=#k��k]X`h{������D$A������dLu<"X�����+\�yy������ʄL]����û��������������$����������]d��������������������������Ɉf����`5f����������������������������Q8�����廯������û�~������Ќ\/++#���W$n��ap�{z����ƺ���~��ѩ�d$"Xh�hXaSWW$n�y������襔�����կ�������������yD���������%��������������������������m����̰`Fc�������'V�����������������~}i������彽����������k�������۶��S�����N4m��{����������ǔ����~L3
7Zh���hpVNnE=��������꥝���~�û���������������������ѧm,������������������������������ܢ��{C!5f��mV

'����lls�����zffudk@8��������������������������������������y������p��������Ld�~L3<���h����yaWk+=�é���������۝�������������m!-�����������������������������������������ш���VM��ܰ`