�{�}}�v�u|�k�e�m�u��u�t�l�r�x��y�i�e�v��o�g�u�|��}���z�w�p�r�v�g�l�o�x~�j�n�|��x�l�z~�}�{��|�y~�|�x��z�z�y�u��w�w�|}�y�r�m�{w�n�t�t�~{�w�~�{����~�~�z�s�p�|v�q�v�|�p�p�x�r�o�t�~�|~�~�}�|~�~�}{�w�v��s�o�y�w�n�u}�u�v�x��}��w�x~�o�q�z��t�u��x�z�z��}�~~�}�y��w�|��~��}~�s�{|�y�{�~��}�y�s�x|��z�|�~�v�{}��|��{��~�x�w�|�|��z�}��t�w��|�y��{�|��{�{��}�~�~~��|�y�y�y��z�|��z�{��u�t�~{�x�{�}���}~�~��w�x��{��x�}{�|�|�|�{�~�}�|�~�~�|�~~�~|�|���}�y�z��~�|�{�{�w�{�~~�v�}�~|�{�}��x�|�}~���{�}z�}��|��}��~�x�|�|�x�}�z�|�x�u�z��w�z��}��y�s�z�~�}�}�}��~�~|�~~�y�}�}�{��{�z�}�����|�{��|�z���z�����|���|~|z|wz{w�v�|����~�|}~z{yy}{~������������������������~�~�~�����|�~���}��|�z��|�|���}�}}�~||�z�z~z�z}~{|~}~~}~}~||~|~}~}~��~}~~�~���~��������������������������������������|����|����~�~�������}}~~��~~�~~}�~~~~�~�}��}~���~�~�~���~��~��~�������~�����������������������������������~~~�����������~�������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                RIFF��  WAVEfmt      +  +      data��  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������~~~~~~~~~~~~~~~~~~~~~~~~~~��������������������������������������������~~}}|{{zzzzzzzzzzzzzzzzzzzzzz{{{{|||}}}}}~}~~~��������������������{xspnoppsvwwxyyz{}|}}|{zywvwwxy{|}~������������~}|||||||}}}~�������������������������������������������������������������~~~~~~~~~~���������������������������������������������������������~~~}}~~~~~~~}~~~~~}~}}}}}||}}}}~~��������������������������������������~}}~����������������}zwutrpooooppqrstuvwwxxxxxxxxxxxxxxxyz{|}~�������������������������}wpjea_]\]_adfjnrvy|~~|zzyxxxyyyyz{}~����������~}}~���������������~{yxxwwwxyz{|}}}~��~}|{zzyxxxxyzzz{|||||�����������ķ����zqmaUPNNLNV^finv{{z}~~|||zwromkihkoruz~��������������~{wussrqqqrsuy|~~|zyxwvtrponnprtwz|}������������������µ���zmbYRLJKMRXajqx}�����|wrnhecbdfjmquy~���������}~���������}|{yxwuttsrqqpoppppppopqqqpsxzz|�����������������ĸ���yj[OEBJPRX_gr{�����~~yrkd^Z[]_ceipy����������|wty��{y{~���yvw}�zsooprvqmkkottqopqrtuxxvw}�z����������������ǽ����gYPLNMIHNboy~~�����skkgbZUV[cgjqw}���������yus}��ss~���}x{}ynkqtrnjinqpoomovzsnrw{||}~~������������������ǹ��oe[VPIECM_jpry������{ysj`XWY]]]alv}������������trz��zstxzzysoswvqlloqokjknqsqosxyxy}�����������������������ο��~s^ZTE<AMU]djy��������ypd^\[VTW[dosy������������wx|{uonpprtqptzzursuuqokkkoonmrvxz|{}�������������������������ư��oomS98GFLQQany��������uqlg]YUQY_cjpy�������������zsjhfefhikptwzzz||{wtqrqqrpptyz{~����������������������������˲����y]NNGHHDJRYcqwv������{trka^\_dcbjsx~�����������{vohgkkllkpuxy{{||{}~}}|���������������������������}����������������wpgiibba_`fjjmlquvuvuruttqqopqrttwxz|}}����~~~|}|{{{{|}|}~~~���������������������������������������������������������������������~|{zxwvvuttstssststttuvuuwwxyzz{||}}~~~~~~~~~~~���������������������������������������������������������~}|||{|}}~��������������~}}}}}}|||{yzzyyyyzzz{|||~~~}}~}|{{{{{{{|||~�������������~������������������������������������}{yxxxyyyz||}~~��}|}|{|{{z{z{z{|}~~����������}}~~~}}���������������}||{z{|}}~�����~}{{{{{}~���������������������~��}{{zxvuuttuvwyz|����������~}|{zzzzzzzzzzzzzzzzyyz|}�����������������������������~~}}||{{z{{||{||}��������������}|zzxwwwwvvvuuuuvwxz||}��������������������������~|zxwwusrssrrrssrsuvwxz{{|}����������������~|ywusrrrsuy~��������������������}ytpmligfghhiknpqtxz{}��������������������~}||}}~�����������}|zyxwvvvvvvvvvvwwxxxyyzzz{{}�����������������������wnifc]YZZYXZ^abekpsv{�����������������}{xwwwwvwyz|~����������~|yvtsqpoooonopqqrrssux{�������������Ļ�����|xna[XVOILPONQY]^dlty|�����������������}|ywuttstuvxyz|~���~}zxwusqpnmkjiiihijjlpuz��������������ô����zth[VTOHCGKJLSZ^_gpv|����������������}{xvvvvuuwxvw{||{||yvutspmmmjgfgfddefgimrx�������������ȹ����{uj\XVPIDEHHJRY^ahpty������������������}xvxwvwz|yxyzzxy{zvtspkjjgedddbabbcfmsw}�������������ʾ�����xl_ZYSLHHGGIPW\biptx������������������|zzxwz{{{|}zwwvtrrqmjigd`_`^]^_befjqw��������������Ⱦ����}qc\ZTMIFCBDJPU_glqv}�������������������}{yyyzzzzwutqmkkifeda^[[ZYY[`ehnv}��������������ſ����vg^ZSLHE@>AEKPZciou|��������������������}zwvutuuurpolifecb`__]ZYXY[^gos{���������������Ļ���ob\UKGD@<=BEJS\ahqy~�������������������zwtqommlkigda_]\YZ[ZYYZ[]dls{���������������ǿ����zi`[PFEB<;?CFKU\bjs{��������������������{xtpligdb_]\YWWSLIIGJACXl}������������˴��~m]\XLKMOS_mx�������ypnogac`[_hpz�����������ujfaZ[^\[\[[]Y\_\]ecait����������Ľ����xpnqhenkmuw�������{lcd^[^dgkv~�������������}yqiiknrtuurlhhebb_XRKGISe}����������ά��tkryzwvpjkkz������}xmfjgc`[\bjx�������������xjdbbjtyxvqhceikig_RICBQg~���������ѷ�{skw���umadgu���������xsj[SNWfq�������������|phhijjnnjmqooooha^YOFCGTn���������Կ�|zo|���si_faj���������qeYPJXls�������������~sdfibcjljlonkklj_XSD8ATh����������Ȋv|sy���vi\a^c����������qdYOGUlu�������������sfffacijjnnljgd`YTJA>I[v���������Ӱ}{w����nb]b\p���������zi]TKLbry�������������xkeecdffijihieb`ZPD@CJ`���������͔yw����~j]_``~���������ucXOHSlu~������������~tjgfddeghgfghca^UEBEG[|���������Ш~z�����o^^c^r���������~gZTLPgv|������������zwmfffcbegedghd]UF<?HWp������������{�����xaXcag����������nZRPM_v}�����������}ysiefb_`gjiijcZVQA<FQ_x���������ǡ~�������i\^edu���������v^RPPZq}~����������|ypeaa``fkiefe`\VK??ERk���������ȭ�������q]\dal��������}_PORYn~�~}|}���������~tf][_fiprjba`]YSD9:Ic|�����������u������y\Tgid{�{������eKKVZj�|wy����������~kVSXblx{sg]]\]aYE;;Cb���������ɴ��������rXXccm���������yZKPXar}~yv|�����������uaTW_gourib`fgd`P63@Or��������Ȼ�~������w\Wbdhx~{������}_LOZcoyyut{�����������xcSS`jqwphggimke_P95<Gh��������ɹ��������s]Yabhwzy������x[NU^dmtsrw������������wbVUcmlppkjoqnga^VH=<GZz�������»��������{f_iiagqy������|hWYab`dlu}�����������odaabhoopvtpmkha\]R<5>Rx�������þ��������~h^ilegqz������}m\Z`a]]hw�����}�������ytfadbbnzyzvpligfaZN9/?Y~�������ĳ��������ykkrk``m}�������se]ZURZn���������������xk__bamztwxqnni`VQI74Ko�������Ʒ��~������utvj__jx��������l]VROUgx��������������}omlia_jux��}rnlib\WK92Fl�������ɵ��~�{���~�k]`nvy�������sc\VNP`ms�����������~��vusihkfitw{��zrngd[QH=3K}�������°�wxrjp������qgnoil�������yofUFK[dn��������~uusuzsu|ynpsjiqzzwzysihd\M?5Br�������ѽ�{of]d|�|����}zrhhu��������zhWSWWYfz��������|wnbfljo}|z{yvtspstrpnrlf_SE;S�����������ucT`pmo~������tqvsns������znhdZW`ny��������~xlgb\\oyty��}zwoioniadg`SERm��������Ү��ta]ga\m��������~ynmu||w��~yvnggknow���������yqb_bimho~���{sqg_agcTLJXm���������¥�jX\cZ]o��������}oqruqpxz|z|zsqrurry����������nfjwiYcrz|�}~�~mdhl\SNNOYn~��������в��q`W]UN^u���������{xwrjbhotqrwx{||{z}����������}ouwjafqpuu}~}vnqf^WWTPNUq~������������}j][NAOeoq{���������zk`ceb]`lqty�������������vpwqkothl{�}uz��rong`YZTRQ\aj~���������˰��{bXOCFR\dl~���������{mg_[TQY_ejs}�����������{pmupjprpt~�~y~�~soph_][ZVTX\eo|����������ɵ���hWLGDGRZfv����������ynaYQMKOW]gs�����������}|pilmegqrrv��}��}uspga^]\USX\alt~����������ۼ����^ZPBAHRUbeu����������|jb^WKHNT_div������������xonpjbafnsvsvyz{}}upjhihcacbdjrx~�������������Ļ�����zrg^URTPRZafiqw~�����������|ywtrrsstuvwz|~����������~}}}{yxvuttsrrrsuuwz{{}~~~~~~~��������������������������{wsoljhgfeeeeefghikloqsux{}��������������������~|yvsqommllllnoqrtvwxz{}~��������������������������������~{xurpmkihfeeddeeghjlnqsvxz}���������������������}zwtronlkjjjklmoqsuwz|~��������������������������������|yuromkjihgggggghiklmoqstvy{}���������������������}zxusqonmmllmnoprtvxz|~����������������������������������~{xuspnmlkjiiiiiijklmoprsuwy{}���������������������~{xvtrponnmnnoprsuwxz|~�������������������������������������~{ywtrqonmllkkkjkklmnopqstvxz{}���������������������~|zxvtrqppoppqrsuvxy{}���������������������������������������}zxvtsqponmlkkkkkklmnoprsuwyz|~����������������������~|ywvtsrqppqqrsuvxy{}~����������������������������������������}{ywusrqonnmllkklllmnopqrtvxy{}����������������������~|zxvusrrqqqrstuwxz{}~������������������������������������������~|zxvtsrqponmmlllmmmnopqrtvwyz|~����������������������~|zywvutssssttuwxy{|~�������������������������������������������~|zxvtsrqpponnmmmmnnopqrstvwxz|~���������������������~|zyxwvuuuuuvvwxy{|}~��������������������������������������������~}{ywvtsrqpponnmmmnnoppqrsuvxy{}~�����������������������~|{zxwvvuuuuvvwxyz{}~��������������������������������������������~}{ywvutsrqpponnnnnoopqrstuwxz|}�����������������������~|{zyxwvvvvvwxxyz{|}���������������������������������������������~|zxwvutsrqpponnnooopqrstuvxy{|~������������������������~}|zyxxwwvvwwxxyz{|}~����������������������������������������������}{zxwuutsrqppooooppqqrstuvwyz|}�������������������������~}|{zyxxwwwwxxyyz{{|}~�����������������������������������������������~|{yxvuutsrqqppppppqrrstuvwxz{}~������������������������~}|{zyyxxxwxxyyzz{|}~������������������������������������������������~}{zxwvutssrqqqqpqqrrstuuvxyz{}~�������������������������~|{{zyyxxxxxxyyz{{|}~�������������������������������������������������}|zyxwvuttssrrrqrrrstuvvwxyz|}~�������������������������~}|{zyyyxxxxyyzz{||}~�����������������������������������������������~}{zyxwvutttsssssssttuvwxyz{|}~������������������������~}|{zzyyyxyyyzzz{|}��zz�����������~||}��soqv|����������������������}zwtssstuttssstvxz}�������}{{|zxwwwxyxxxzx��}}{vstpopnkghjkostuy}�������������������}umcYROPU\cginu|�������}xwvsojgffjnt�����������|od^]_ceec^[_hqsqrssvz{~��{yxyyz���������������ÿ����~k]VQNNOOPWbku����������}tkc[XX[`jx�����������wi^ZWUWWVRRVY`hoswy{}�|xx}�}sim}�������������ï��seWI;23<GPWamz���������sjbZQHFJS`p�����������xdVQQQPMJILSX^hv~}vry���rnx�������������ɺ��|k^QE:7;BLU_kx����������zph^TLHJQZi{����������~l^VTRLFDGLT\adkqvx��|z���������������̹�yggjaQC<>FVfpv}���������}zvm^NGMYhw����������}xsk^RLKMRUTQPXforrpns����������ͺ���ʮ�{qmniYG>DTeszwv�����������iRJOW\dpy{����������o\QQSNIHHGIR]a^]co}�������������к�|ple^TG@FZnx}�����������tg\OEHQYaq���������~riaYPIEEEGKLKNXcgefs������������ç�}fVQSPD?Ke�����������yqbMADLSU\p������í�{qWFOXH4=PSMKNQXbf_as�����������¨��hXSLC=DUiy�����������ubOFILKLWh}������ƞzlTOTH:BUYQMNS\\WX^hu����������ж��k_SHB?HUgy�����������j[OHIHJOYl������Ƹ��ygXRIBDNVTQRT]\RQ_fkq���������ڴ��znQD?;NZalw���������~naVRH@EO\gt����������mZTNEAGOQPRSVYV[eci{���������é��{^LKDJPP\n�����������|iZPLLMPR\t�����ó���|hXOGFIFAIVWLLVbegkz���˻���б���sXTOOMCH]u������������mb_[RHFP^iz����������sifXKECCJQMFJX^\`hw���̳���Ӽ�Ħ�ki`SM@CUemlt����������~xjXLIQUOQh������������p^SRMB?FMNLKOWeldp���ı������ɮ�usk\N?BS][Zi������������vbZXXPFI[q�z���������xnaVKDINGDMVQRYflmz��ô�������ä��}i[KAIQOKUn������������ynibUJJPX[i|�����������~m\XRJGIIJQPQU\ehkx�����������ͯ���t^RIHJFDMapty�����������yj\RQSQNWe~������������|gXUQJKIINWXTZfkiju�����������м����h\WOHCAJU`fp�����������uga\UQOS]ep�������������n^]YNLQOPY_\]flghquz�����������ɽ����oaWNJFEJT]gr}�����������vme_XWVY_fn}������������{l_^[TTVUX_eabkrhhptpz����ï���˼�͵���za\VLGKJMXgrr�����������~rkhc^]]bhmv�������������tgedZW[ZX]eccfomemuni|�����á��ۼ��ȧ���n^\QGKNEO_olo�����������zpmjd__^fjmn��|��������}�yfchZX]\U`fe_gsleqwolw�������������������n^WOJLIKV`nnx�����������vnlic^`cijpw����������{�wf`f\W[\W_gdblskirtqot�����ȷ������ɺ���}eYWOJLJRZdpp~����������zqmmhbcdhmps��z�������wx�}^^k_M]_UWic`dvjilxnps�������Ѹ���ï�ƣz��lMWXNGPV[aswx�����������qjnoechnoqw���y�������o~�fXddNTbXOei`^nthfvxkt�������ý���»�����zbTRPNMPX^iuw}����������{olplfglmqt{�����������}{thc`[WXYXZaebgnngmtomw}�����ͺ������ư���o\XRJJPQX[qxu����������wnmnigikms{������������}vnfa\ZVVYZ]bcfkmjlooosz�����̺������ǳ���o`YUHJQSWYn{t����������wpmmghillv������������~woi`\XYVUX_aacikkhmpor}����ƽ������˻���vc\WKFPQVVfzu|����������xrongfhmox}�����������|tkf_]ZWVX[^`acfgeiopvz������������é��}k^VPHKPTZ^vw{����������}tqnjfgmtvx����������|xtlb_^]WXY]_`abcefiouz�����������;���vk]SKFNQSYewx�����������zsqojhjswz|���������}uqne`]\ZZ[]^`ab`afmou������������ĳ��{pcXNBHNOW^lu|�����������xtqlkmsvx}���������zsoke_][YZ]^]__``chko{�����������Ǽ���wgZQFHFHQZdlr����������{xtqrvwz~��������yupkfcb_^_`abcdccehlrz�����������Ƚ����xjaZVTTVZ^diosx|�����������������������}zxtqnkgeccbbccccddbcfjox�����������ƾ�����wnf`^ZWWWXZ]`cfnsw}�������������������{wqmjfcbb`_abbbcca_`adks������������������yogd^WTTSQTYZ^dntx��������������������~zupmjgeecaabb`ab`^\\]_gq�����������þ����zofd\URQPNRWX\bmsy�������������������|wqmjeaa`_^^]\\[YVUSQW`hw�����������������|lbaXNHIF@HPSS[lrx�����������������wnkhc^[WSTUTSRPLJLLJO]gp�������������Ȼ���teZVI@?@=;ENRXft{������������������tke`\YWRQPQPRRPMNNLMPSax�������������ɽ���sh]WPKB@@BFJQX^ju������������������yne^]ZXSNLNSSUUTRQSTUU]l{�������������ų��}od`XQMIEAHMPT[elv������������������{rica`]YTQRUWYYYXXXZ\[XYj�������������λ���vmaXWXOFDIIIQXZ_hv�����������������yrlfcb`[XVWW[]\\\]^^_`_]`�������������ο���zufa]ZNEJPONRXW^gt|����������������}xtokgea^[]\[]__^`bcbcca`e�������������������shb^[OKMPPPVXX]equ}����������������}xvvsmjgeddcccccdghihijihiv��������������ƻ����wngc\TTWWWY\]^bjmrwy}�������������{yvuwvusrqspsqomklmmklklnnqnrv����������Ŀ�������yrmhb^]_aegjkopvxz{{z}{|||zzz|{|{}{��������z~syqupsmnmopts�v�{~~~}�����������������������|wrmojnmomqquwyzx{x|x|x|v{y{zzz{{~~~~���}|z{xyvyxvyt{s{y~|}�}�~�}������������������������~zxuvvtwsuvuyx{vzvywxuysxtzt{x{{}{�|�������~�~�{zy}w~v~t~u||w}|�~��~�x�z�z�}�����������������������}�wywyq{mxrvwwuxxx{x}w}v~wy|~w�{~{~|}|�y�x�}��}|}�~}~w�t�z{|~}�}{�w�x�}�����u�u������������������������}yzvvwyvvqyyw|x{vv~xywztyyxtz{x}~}z}���~�~��z�z}�|}}s}}z�}x}~|��v�}����|��}~|����������������������ztnqqnrnoqmxvwuxwx{{|xs�r}|v|yv�}z�{���}�~��{�{}�||}{uy|t�r{{v�v{{x}||��x�|��y�}z�}������������������xosifja`hhnnpvyy}�~}z}ywuttpswuvzy���������|{wvvrrwuovuv~yy~yz�z{�y{�|}�y��z}�ru{s��������ÿ�������mldjeXWc]Zrqqsx�����z{~tojmlhlwpu|�����������~||suqnmlptvrww|���}���}||}~~}~���}��}�|~�}����������������{w]YbbeXZ^njw~yz����|~yxwunijntxr}}�����������{yyormcirllvst|z}�{��������~{��~��~��������������������������{wumbgeka`hxprx�|���u}}�tsptuszvtz����������|~zqlphempfksswy~�����|�����|��y��u~�������������������������������|wzrksvnkmuurv{xw}�z|��z~~y|z~�yz����������x~}zsmlojipmiowzyv}�}���������������������������������������yxsvqononmqxsswz{z||{{}|}xy|yxzyy|{~~|~�����������{xuopmfikhjmnorwzyy~���������������|������������������|somjecdfiiijkloprtvw|~�����~~}{zyzzz{|~������������~|yvsqnljjihijklnqsuy}�����������������������������������xpgc_[XVURRTWZ_ejpv|����������������������������}ywtpmkjihhhhijjklnoquxz|�����������������������ǲ������{qdc]YUQOIKNORYadjs|����������������������������~zwrmkigdddeefhhhikmnquy}������������������������Һ������tdb\VQJIBCGGLQ[`fpx~����������������~���������~wtqmjgfdbcdddfhghimorw{�������������������������и������|rbb[SOFG?ADCJOZ]eow~|�������������������������}ysqmjfedaabccdfffhloptz���������������������������Ժ������~pa]\ONEEA=DCIMW_bov~~������������������������}|wqnmjeccb__bccdeffhmqty~��������������������������ǹ������uf\\ULGBB=?BFKPZ`jsy������������������������~|zvpmkiebba__abbcdfgiosvz�������������������������˽������ui^\XOJEDBABGNQXaisx}�������������������������|wspmgegk\XjbR]f]Zajddx{q|���������������������˾����skgVNHLLHCGTOQZahmw|����������~|wtvuvwy{�����������~wqlia]^ZXY[Z_badjnosz}���������������������������{ilZMJIHDOLIV_^anry�����������~xuvtqpstwz{�����������|tmif_WXYWW[]]bhijntx{z|����������ũ��������į���p_^TLEIDHVQXbgls}~��������~xtvrppmotuw|�������������zsia`[UWWTV\bbeikpuxwvy~�}zz~�����ƫ�������ƾ���y\WWK?BKIU[Zityw��������ywtphkpklorw{�������������{ojd^^\QQY]\]cehooquwuv{zxxvsy�����Ǻ������»���~hOLNJBGMO`gly���������|xrlhgd`gmnqu|��������������~yma\Y]`\ZY[^bkmlkjlqtvsrqnov~�������������¬��wtgPGJJGPafotw�������|ywrjc^\]`aisvz��������������{utpjc][agghgebcikljfefhjmoollz������������Ǯ��kbc]NISWT^p{����������rheb\Z\]adgp}���������������ysqqpnlifinpqpnidcbcecbbbadhmo{����������ž����dVTRKObjfmz��������z{sjbbaXTX]dmt~�����������}����}zxutuwyututqnlkhgfdc_[Z]aceikt���������Ծ�����iWROJLbwy{���������|um_WX`a]`ehkr|����������zx{zyzz~�����}vuusqolhecbdhiihfb__`dq����������Ƴ���{l\WUSS]p{����������~wqg]WY]]aipux~���������}yvuxz}}|~}}�}zvqmjgdegggjlkkjfca`an����������ï���yh]XRPTap|����������{wpf^YXY\cksz~�����������}zxz}}zxxvtux{}}{wrlebacfilmje`\ZZ`p����������Ų��~qbXTPPVbq|���������|vrld]YWWYakt}�������������}|{xtrqqqstw{|{zwrkfcbaabdd`^___et����������í��zn`WSMLR]lz���������yrnia[VTSU]ht���������������}wrmjijmptx|}|zwrmjgda`^[[]`bchr����������ϻ���ui]XQKKPZds���������~wqh`[VROQW`ly��������������zrjc_^`ekqwz{zxusrpnkgb^]\\^bhr����������Ƶ���sf_UMJKOS^ly����������vph`YVUUY_hq{�������������vld_\[]bglostvwxyyywtrpnlkkknt{����������º�����sia[WSTX]bipw}�����������|wsomkklnpruxz}���������ytrrrstsrrrsuwxz{|}}~~~~}}|{zyz{������������������������|yvtrqpnmllkkllmnnopqrtuwyz|~�������������������}{ywutrqqppooppqrstuvwx{~���������������������������|yvspmjhfedddddefghjloqtwz}����������������������}zwtromlkkjjkllnoqsuvxz|~����������������������������~{wtqnkhfdcccccdefgijlortwz}����������������������~{xurpnlkkjjjklmoqsuwy{|~�����������������������������}yvspmkhfeddddeeffghjlnqsvy|~����������������������{xurpnmlkkkkklmoqsvxz|~���������������������������������~{wtqoljhgfeeefffghijkmortwy{~�����������������������}zwtrponmllllmnoqsuxz|~������������������������������������}zwuspnlkjihhhhhhiijklnprtvxz|~�����������������������~{xvtrqppoooopqrtvxz{}���������������������������������������}{xvtrpnmlkjiiiiiijjklmoqsuwy{}~������������������������~{ywvtsrrqqqrrstvwyz|~������������������������������������������|zxvtrpomlkjjiiiiijjklmoqsuwxz|~�������������������������~|zywvuuttttuuvwxy{|}�����������������������������������������������}{ywvtrqonmlkkjjjkkllmopqsuvxz|}���������������������������~}{zyxwwwvvwwwxyz{|}~���������������������������������������������������~|zy