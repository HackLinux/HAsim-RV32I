������U3K���ܬ�lV��e�(Gr���a�tM�ldks��hu�p\cr�������m=�p_5��o�NNw�Mzw����!hS����8q�Xa�~`iJ�3ò�S\��z6�|c��IMȅ��=!\��p�Ǜ1�ڐD���C�F�W1Q��Fɷ��酱	n(��v$c�<oiI*���1�2F�[��D��2�v�$��k�\o�Ռp�@V9��c������~�n~��h"���[G:�`yn�ZC�Lq��ff_��m���W,Y�r'��b?Ÿچ�P,wbDn�s2�Y��ZqKZa�Z��[��m�!d.���*)6L�hz�/0 �\�6M�^��lȡ��B�x(����(���$�1p��![�LQ�qa�� �5��W�vd���
nᬁ݌»������s�3�GY�a�&v~�����������2�$�u��k��ѐb1�N<N������&���F�M�F��N��}�\k��~�f��n�unw�j�:h|�XNQ[�7�b�V�b��5H��D�oBQ�xa�����D��Pan�D���m�k�ڙ��6�j�v��h�"S�N|<�y�J�2)�u������`ge��X�RN�����Έ�u���M(����t�T!�U�a���+a:����M�K�P$2iT�b)\V{A�h�d0��������3nEy��d5��Ť|
o�PmFo1����pTI9�F6�5S@�p�k�-��$�D��"��[�}8o�2���&E:������|�|�5���m=}�κH���L�˫�0ц���AF!�9��*i��Z���jl�hF[s������ϫ��$�H��-�o�r)�q��6��K�ގs������V7j�Opǻ�w>ж+PJ�:�OQ���-�>|�w<�X9~�����������<�?�굄�q~N�@�ހ,EߞF�(dw_>A�T�H(24C�8�՞M'���g��4I��<�E��Y �m���>�|��$�r]�YO!���w!�����	i�Z���=�0�B`���wx�����p?�,{[���!|�����4�a�h[C��Ed]qw����zu/\FY`	�x�7��ޮ!�K��/�c'a�Ʋ����	yyZt@~�����M�i��x'�&�k�� ۥ���Ʌ�"d���}P�O::�s����4$�=�/�#-�q%2�M�9<BZ��X}o��_Θ�po��+-%�j�k ��Hh%0f�?�q��JjZ�%����Ȍ�'��)������<��Rײ�T:�%)w�V>:~�as�	�gO�O�8��yN�*��a."·0W.&`��ߨ�2�6��v/�R&�&w�9�^[S-�:�����9���8���ќ�<y�����
y����[)�Z�GK|�[r+~ |�H��F��*��]�+��E)�|�,�����U`�H�(��=�Q.G=|k'e�O���`��̠R��s��&�_<�ߖ���B�l�HҲ���=Q�t�0�%e\�G�\���>$iN:R)s^�Z+(�����&w���t���?/�Ͷ$lQ
ߤ×v��h��V�ϐ(��5�lN���S|
��:3��~�~K�cT���-E�vS���N��=�w;��f7v�+�G*nhݻ�+<���ĵ㛹}�Tʥ�+�6
1�ѾBV���������h�����wط����8ђ�kk �r�������%��$v��;���4ؒ�k����S�Vÿo�'N߽�>�� bKD�gF�*��� �/��`3%���e�j?;gO�����p�b�Q�Җi��^},�Z&�Yɂ^q
�%QD�w��&#[�eI��&G�kL�V�W�ڬ��*lw�,i8Q�I,2��+�#��U(�P���)�1�a���5}!����{�ʠ;�M���g��{zp/��z�W!%Qn_��(���ˮ@���	cFn�q��6)�;�s_[س���o{ş��_t��_�z�#���m�j����4���BrZ%Y�inܨ1&ǩE���Nڌ�l�	�խ�z�	T��˳�~���!c�O<*��0çE?}������)/���i|����9���8P�ݏMڴ!f�ޣ7�����5H����_�B6,<#	O�ɞ/Њ�ي�B�B�X�I�p'ܒ'9��A\��Z�4މ�k���꯭�/��������[���W���\�}���z2��|�3�ϑN���"��c?����@a�_�8KD��!�=��K5�	Q�0IX����q�zĠ�Jj<��#I��	�#H[�(����j��Jc���85�l���y�FH�q�������I�eT�n���jj5��A�/�%�3B;=�5haң�����%�,��2��������n$9��#�V��ÙV"���jC@;��/!�e?��U��|���L�S�K�F&�U�q���T�k��K4���E�!d�|c��/��j"�pCq���D��"�j����)��AnVf���6A�Tېx�7t��7�-�-��`�[2gJ��SG�����vof-z�a����`��8v��%�F(G.�2��ɕ��u�р�2���1E�N= ���P��g	=O6[n`ٷ���@�4d�Ƴ�����)��ڡ��솻Mȕ����ɲ|yp�Чc��%kP�@���� �w�f*��?����z�F�YM��ArcBѦ��`k�hS�{~a#KU��ƶ����7��O��D�]�ֲu������muc�3�<�u���L���%4WM�{��*``�33��b�N�Y�Cl,���ɜ�&G�i��~N�1��.0wV��,�b�c�Af7ī�T��x��E�?�����8md(Xæ�������}\g�W�q��j�7b�������/&�OZ;���O�r����	&L����PYBU1ۊ�0U��R�sA�A���,W�����}�y=���zl�<T���<��O�"߼<��.8�'�r��X�{#�k��v�e;�G�1"pu�N��@)�|�p?�nfkK���/�uecn�~���� �縒=�u�_����#��,b�AH�o����ҨM<��y�ER3Zs<Wė>�5�(*�4{ۥ�����?���w)N�� �%�-X�}mc�=��M�t�tW N�럏ix>C{��ƿW�R�f��'!9�Rѽd`S0�,eg�F�_C�rL ߔ�oqֿ*�$�9Q��Aߑ6��Y
�����8}��/lu�NYJ����p�cM<�b�u��.�no>��:ہ�w3A�����֕�Ө�w;�/��ʹԴԑq[�uf�B�R�D�'"A���$�! ��A�$�M"H�".���]W鹲��F�����Ry�R�V��㩣U��c������:i'��0��u�ӿ�v7.��!������b9=�;1��@!����xn����F�v���d`����s���.$�P��p�v+�6��V���x ��Y|�(��c�N��uOh���w��k��֩�{� �=t���{�uUr�O���������ø�������]^������ {�?�DfJ��<*$wU��L�!�pv���22��������|�֋�´��(�ym7�PX��~;{��H�����6��|9:���������0t��v��}��;����χ��{�tq;���}9,��]�t5߱��Tu?��s�su���ڢ���&��y�i�j����5&������z��׆���c��뵵
�7�^[��}r��=n����9��_�w���������wu��r�5��p��(�%����-��sঽ��
�䋣�+���y�U��H����|f�y8��:/�u�z|���E��5_3�V��#�-��}/�H���9V��
�xS3�f�{Hǰ[�6נԖ�w�$�w�k^߭���p�M ���8Bծ��z�{������[��u}����J��#�T/��*�E��}4�vL���z4������nu��4i��v ���~��	G���b>��xq���A��>�ٚr=m��i�pț�1��Zm��pѫ���p�_�u?~���;���a�nW��ؐ��݁$�v�����|���͓y?��>���P�)��A|��}#�A��������A~[���� ���B|��!�� ����܅y{�	����A~G����m�������P�An������7��C|�����f�롾��A}���C�)쫁����3-ֵM<���Gq��������F}������6	����`��W��1ކ���x��&���?�
�Cy�G{���'��藃��Ez/��ٟ��(�=�Q�:���@s��3�О�;�㧻�m���\�AE�򓛨Gf1�[�ۮ���f�א��D�7]7ҙHb�9����p��5xw�T;� ��!�5�P;�~������8Ĕ�b��;�t�B��K#��d|�y�X��uHI�`�.�@�;��I���z�$���Dzc#7�a�Bvj�f�P����`�Vα�bY���5M�3:�9��N̢= �H?�}�B�h�)bnI-�F��|F2���;��k�/�l m�A��'5��{�5��:�Ӻ�j��]����{��Py���� �[d}:�P����M��*����ua�f=�E�:u�7�A�k3ő}��Q=�4T�D3�Yk�>�7���$IiM��!į�;�=��>��^�R�?R�f�~�:u}.�=�M��������L���
3�|�̺IFL�t��ƾJua/�Gj\�LjJH���^������������n�|����"m�]M����"-��()���K����:�LIʽ�UN��Xl��ۙ{�c��]h����p�x$� L: ��[h�.�!ܟ�#�p����L�>V��0s�!-�<]#D���E
�b�)�Z!w'A��u�ڜu�+��mގ:�W.I���;	��a��=U���{\�a���)��B���u�����iV��"$�1���~�,1��(�\��%֩���XFư�?}�Oq`����_>C��T�Bq�Y3yZ1�|�y�L�r��?�Z:�0�P�x�E��\��ǻ��A�p��"��������^5�l�32A�G��3g�I�I�_�!�����ܘI�ag��_�Me�1���	�q���	4K�q�쏕��'��j{�s����"�ۖ=qt��_��v.1�{{�P���f^��/��z����E�Q��� z��]j�\����� ��	�_�i[��Op1&\ٰ��u��L�=
�C4�~ �y�B%�Z���F[�<p�0�����{�RYŕ}�Hk�qΘ��&�EL2ڸ�|����=�lt�7K<F��$�dծs�� 7xR4X��N,�����D?4w�ذ��i�K|�Z�D�yN��gčۓ̒���B��ty�7�ܙg�Aܥ/�̒|�	���X>���ӂ��'hy�`5,�mDvK:D8��0��خTC{���7tc��D�>����E��@�,s1+~a�Er2���s��8[wco⨰R6��0���.P�b8����e���AWVK.�}�C�Y�~�?gXr�{q-���ku}[��QY�{��7K�\[1�@5؉�0:���m�d�x�:���.�Q�������8W.���(f(s\�-11��%��_���V����e����F"�D ���u �Vg����$r����E�eB#mE��m�@Sg���$N�42'@�:����^����{5��<��>�l�n�[\���4e�l�ל�&#���A�m߀�rH-�vKUQ�:�]�q����tlD��~b�薚i��Toc�ìm	|�>��(���A�w�2��𚩙qﯸ�R~?/&���/J(��zNvj�]\����]}�۳N�������X�ʉj�޴*V����R����Y��jTyǺ	Gf�^ 6=* q��q�n�V=e�az,Ik\ +��I}��ݓ���Q#Ơ���QH6M�~��i���%�L�n\cU&��͐rW��S~&� �����kCy6d����_�t�����e��ަ�1��D?�x��"1rQOz/ҐypO��h"ۙ������	�Ԇ�Y�q�c4�JX�L���.�C�8�~ ������/j3]��@��2b�x�P����P&�I��`�����}��V�3�T��Z9ɴ�M�Q���.* �z�a�|8$�]�.?����ԥ����\n�J���.mk�א�fڝL/��U\C�5����Ì�Wiy���^���r��=�8�����������/�v�Yyi C��0����=r3���Xy��|yy�����3�.������<�K����j�}��{!���ؿ(�䥻���c��&鳐���:�Cz���{.�y������άA0����ĿI�o�k�vi礱}���YX���5�=}=�9\����B���k��!:8l0�v�����|���O��3��%X�4pk���p��#���ߠ�#lE�^C��%Z�5h4�]���T*i*D
�c��2<�����D�'Bӗ�5�Ƣ�7�C3�[�[�Ӟ(��R�:7�6�m��+�X�/��c���H���%�#�+�%������٣@����b"�,��e�*�˘����EEƷn{rg͵�+��.����I]������5��|P�a_U����)*#n���(08�OH&d�\�=Ѩ%-����)��]�]��h&W���.��"���A�$����D�v�[	���r�ϴ4N�5K(�5_,�86�j�E���1�����G�WX0��(�GVQ$|��'Y�"}`3��t\hvp-4@�`du��Sh��:ز�=j�TH��!�{ހ+39�ܖU�3��@�����c?%'�]ݭ�z|Ų�еa	����-ɗ�'H���vE�]A��AP�:���8��˻�46�w�Ae�و$y}T��řwvh���J
>�Q�-����¸�}b`�moF�J�hR0?wb���¹)��;u�l�ۑ$S��BV�M�%3^�N[�I�ρkQ��Z�&�aO'�0��G'��5ma��d<ɦ��r�N��\��ubYd��e�҅����A֊�ǳy���3���b~��S�PpBa#4��
�:͕ /?�cw�����~�ZO�.���]r�*�d_~���R�5�W���ӆ��w��S^O�a�:��hh��VG����R�|##$%f�D����U V����Ui�*/nʵ/��d���%N��h�<�|uG�6��*`A���r�����ꣳ��&���vf���Tz���e����4@��0Ͱ3{H����k�_��r�Q���;uf�ɑ�Λ]�ξe�'g^�����]O�gǍ���n�pf��I����pze�r�C�G�|��!��eo�'[��OEO����]�N�G$Gg����Ȋ��njUa�ɵel��,������a�����N��\Je�'��T�(�����_ݷ�#h1rv,�Sg�=��F��_�ۈ�3nd�o�t^D K��hȗFZZf����;i_.�o�l���¢s}�<E���,7����r}|��I�*�����7��#�%�H}&5��M���(IٻilO�����zW�_���%�Zԣ��D<��5��'�X�a�M������bM�w��j��p�l��G.��<ܸ����B�.�]��n�,�l��ښU)�c=�x]3٣\��9?K��x�c�@%������b6�pF.^ʓ��%W�f��TК]�._܁��.|A!}˷��=ǉ%�qJo�o�����»S/���-tim�ر�P�G�إ�(��W�����_g�̴���AV��/#fb_���3����K��I�Ҽ�I;|Q�4Z�b�2*	E���,�އ�O<�(�a]����ۚ����^l+�5\��]iI�]�;�R�hh���Vq�Vq���h�,���r7�]�d�&��6l�Nh�k�T�D^ï�$�ےh�����D�_�����R�D@V��c�g��jv�?��:�Y����Q-t9���x(2>���D����B�؂�����_�t�����+]�;���=�2��}� h��b-L텃�|Rh{�z-���dz)�[R�?���w{Ĩ#�ۿ/��{�igO޶�-
a�	����i/xح#7��)8���)�=�ǥ���e��qtm���d[��ǣjr��G�:K/9�}j����#ٸV=�)�W[-G_@0��졵e�&_��+w��KI%�������7�8m�jB����(�'���3�g��Ud<l�o@�����Y�x���)0�.�|��t�h�>�����QLt7�Q����}���_���� |p��4���E� ?+��fRWpHQ�ƪ��$]!<��˕S@P��w|2|���sn�,�>�5�
�Sb\�Ũ�ob2�Ng΂<�;b!���e2L�T��3�I�	�v�b�M��ơyk���(�|��v��l��ד�q��#ݡ����狜a�'Pxu�kh��-չ⇕5�;�ܱ��'j��- 
E�ݫ��^i�/����_@b����3u�>��,���f��v��廦4��s�K>۱�+�S��k���+ȜQt;�1!/_�'"hO&eF�B�R̵���|�8Ѻ�+��O��U|է}��{�s2�U�C)F��G<�%B��%\��
�YѤE'ҿˏ�]��U���u�r��Ֆ#�5����և\�Ʌ(_�:���_d���E?]j��fF��,,_����ӻi��[�����u�"UG�-�)���1%���/����L{�A@q?�Cg��{d@C\���J���趈��̸u�O�EX�mr�t���v��U[S���Ӎ���V%��n�ptm.i.M:�e�0�%�j�T��J#]w�M��ɀ\.<��l7&�~:�~D˸���!t��`�먻�}��������ܸ$�D�:��o��VS����{=����TA���]?���O6����RC������#�qQ�c&{'��ȸ`�'qe�M�
<ڮ�{u^�~'�ύR�a�+�*+��e�}3'���?��5�k��:�2~�}��*S}���W�aK�+aX�>4�v4��XT���.i�r�#����=�/��/@z��䘹{0����e����R��F�r���0C��輽�=E���]��&�D�������h�x�o{V'�Z8FjO0l�zϖ�t����߁�R�V�~.F_-.�A�]�_H
S[���|-.��v1׵���^�\��^����F�Ny�'��j�'��-��e�F�}w�x��֫ݾ��'�`[��?�wɲ�F`�m��4v�_��{R�<\>��(����t�^*� J���85+Ơ��?�������}Gs�ߍnc�jb^��'1�r�>�vؿp��`�LW���*�����C�&s�j�[�c����C|��,�W��?��l2�fn��E��,�:��Jc+~�3}��t�3���c� F��N*��������uW4�i��E�ܷ��H�oR���7m����֋��z���ʏ�����$im�x�\щl�T�uݿ-]�__����LPCk̂��-��v��}�y��I|`�
�	"�ԨA�
�e�=F�<��� r#�9�cU�>�/�����f��mkk=l�[�]:��{g ��)k�y����~���y�~�%�K��E�x��|�꺷%`��aS�#�Yh� pq�p��V?�>���a3���e���0y$��K�cz�g9�VTw��Z�P=��x1��\������S�7���VH�n:�V�;�(�:p���U��I�x�{����cس����%�-��;9�W�"�|S|s}�����H��e����!����u��:�Ѫ��~�U�S�u��|?��ш�����xJT���9k�LC�L��մ�"�8s;/����x�Q�vc��lF�KI�����]�X��W�/�z=n�͉��]�,/�=��2k��|����QJ�s&e������Y���R�Zs(�q�����7�-{�����,+���G�����y�S���I�`����tf�mZ�)���8�{n�zIB��p �����nY��$�K�ͮ�zI��|=�ks1O+?SSI^���<{觻�W.o����1T�t��
:����;���?ˑ<�I��V ��EH�T?^t����JqX����=ȍ�ZPw�~���y��Z[�.P;��՞�[��H�-�.�9�:)�aڳ/��x��C���i��@f�����L�t��pi@k;�ڃ��'c��,�I�WY\B�����̜� �M��>Ƴ���dY�������(�W} �"��3�����][����ݽ������XT�m��j�}H��cKq2>��-����cZ����?�m��;K�Z������]BK�B�۵��t����:�\��-�= �a��<_|\�:7�WH!�E>Bq8���b�v[�����񹈁��9`��П٣v ���K9f��njL=���,�/��Ϭ��͓� ��Q׳{��lG��E<T��D3������I?�����=��)v.Ɋ�r:z���վI��xa�u������!�E�U�^��o-��7�0��9ZC�K��۬��⼂S�$�����'�����E�W+��%zy�����3c���;��m����VS�Vg�=�,pۜ����e�	�K� ���XF7�Ѿ�p���$&k%�.'�_�,&���1��j�|g\oqF,��P��q�2l�d�j���9W��Cݏ
>��N;���(v��	��	�S_�.^#�Ʒ��1�X����Gf�&1����0˲�.�`2U+=]bٿ���Z狦��q�y8u�v�V�>��=��(�V������v���?�n�_^��5�/����x)
������q�{S�����"r�	�$�&?�D{ՓkF��K�+��K@�b��*���(�
��N�1���>!��׼N8��yEJI:Ov{|�S�r�#�륆i�bQHW�C޹��IZ'����x�Q|텕�������m��U:��Y��x��!����v����l��<b���uH�ZV�٬Pj�O�![."�Ɏ�@Y��Gu�c(��r�h�.�<�8T
v��Cg�h�;ك"��!�)�l�ڴ�Xw[����������j�˳�`�X���j)�cz�%�&R�y,�%�䜵������o��|��qXkeٮ��������:h���pl��<C~oo�� [ mR�g�T�*��������OE.VЄ��p�����5R�J����U��M���^ɻ
V�hZ;�8�)48����ڿ��S�^$�%�}����fň��4�R�r�I����w�wkTc$6xTc��E�ILۇtW1F36���tQ��y�cS_�a`��E��n/3æ�D8p#��m�U����.�W��)�7����V�x�`�Nzd��<��ꎣ�*���<p�޺��Y����nr��i�cl���4�ji7��M��?tc�}����6t7te�߀��v����F��m�4�)m6E�q�Hْ��ܙ{Q2.��P��L0�جq��F�Yq-�:%�f��I`�y���^��1��LY�w;�e���q�vcuw�p
���r�������n����)�.��X�uk�̎j��4�@4���`�`~U��~��|�Mܒ���A����AeǺ�r��S��h�����yyHZ�J��(8 �3��`����N;�N1�/\�_�Pqi�|�-�����b=?��f=?��j������ ����zw.���궧��Iz�.M��R	%�TbS��H�$-lCvk{�*g����@����(p�ӇV�%C�h��^�n��j��A
��U�P����rw��Z��&�1����-m޶�I�֢(5�˰��t^�ϯٔlQs�r/��sc��&5�X��wb@wҨa������}���t2�J�n���u����c_��A��e�����PS�,�ӮjK��dl�ܮ�5���s�Y*k�@�c�a�wƋO�9���f����@y)��^I��h��t���E�������SK��\h)=؈
[j[�Q��K����ޘ���VS!'��{��o����O@ζ}��a�@P�P빭�pQ��t�
N��ӟ �l�֘���B�7d�����>���s1K�XoT���һ�u�[��Wk�9�����O�1�j�w#� ��;�E�a�����PÄ��~�|_�J��ZA��ٶ�
��h�M�c7�I�jM��j�]�3x�����q���yG�k��q��0uτ9�H�\K��`��~��
z�pk�((�!������ !����!�3"d�'1�ىf�
�5�/�4vĦ]Ў���!Y�D+qMf�gy���9�i�j�<
� 
���gJ�@�T�a��#�����f��}έ1 ���zU���y�D�4�ITb�~l��h�#�;6+�%Wo���`��f�"p4�F�i���|W�ƽ���|ۀvاĿ�բ�EcO���5CsY\Z3B�����0؆�]R��/��4�١E��9�~��6�c�7TC�{�����Ke��宫
�O����jl�-s97V�w-��!�j.+���e�'*<�����%gƋ�E�KI&����pw�Q���a����t�@�9�����G����E��vM�&I�sX��t5N�XxQ�3���խ����9�� �τã�Ͻ���7�'���-�\� 9)q�G���#�9��td���m��}�D�wg�G�b�������}~,L��T��1t��C���,��St�}����c{+�}҄�D��P& �ٙѡ~�b�Y&�K�'�Di�Zո�)���܄�lyq�s����re��j҃��cn���D��ЅA�)6�O��Fyq�x�����h�v��H/j-\C���j��e*Y��O� p1C�����M������fz�L!y֓KB��?1�eψk��}-�o�t�����$L9�x���;���uqy�J�*��N�B_�K��]��	�1KE��
k'�%($?�t���Զ��Aq���me��8J���̼:wYܵ2K0<�I�xp�Y����v��3��g'i�j;>.��#*����F�U_=N����~��L��r��|G����R���N��>��y~u~����N��>~�i��e��n"��5�q��Q���Ӯ�;� ^�\`��,���}iɩ5�����R}�N����-)��k��>�9�}�e�lż}KݞM:Ca�A<��Iu�|�,8�2ȉ혽���(b�`p�C!��}��KA�+���,l�۷���։�8� �Ǿ�T��uFX�k��?z�U>��С��7�'�J�GS��*�xTO
��Y��,3� ������\���EY�����Fe�ꋷ�hR��)�?/���G�$|������&�]q:0��;'H׽�ߨ�G	φ Ί�=�xv�_���oԳ�4����Q׭�[aPRO�rv���lESf�8:\� �}��� �|�1Ԝ0��J|�������qj%,���g���W|F���sq׭:��%�V�]������������I���R��| "����~&e��8vvr�-����r��	q��b;T��}�Q#{)4��ʱ N��4[a2��D{ύ�5�.�K,:�L~b\��,�ĉO�qK�娓Xc�4As��%'�����*GA%���g�Muu�V�`� ��.iwPx9�n���	�����5��
,��5cHA������3���rn�^�6��qD�@����3a !��߂W#��gV�48���*;#vĐ��@!Ď(��۠1ϔm��` ���|3�S��	�8r�3wtx��l�����^�^P���c�hо�
�9�]\H,�	T$ZA�$7�6�)�l��h��v'��F��L��0@6 ��)�7v�P'�� �Z�� ����m�p8P!�f���.uɄ+H��L�}Ċ��H��=�KjF�`M�b��Ϝ�&�j���w�8M�X��a�y�2C
�+�}����J���G4Ni��w5`�,E��d���)�8���$EE/��%��#�Aa�����1Q7i����cJ�k��,���XC�IYh'=���Gr��M�"���Ӊ4�I՟�I��[%�~%]�tY�<��c�'����;��1pK����
�t���Q���	=��D\��X�Mi��h�Fy��wn��Af��Ϗ+ǚ`�<H�R݁�ߗ�}½�F�#���i�eH.zV��[�����17������~7�#E��)B_/�Sm��tWr���qr�Re�х�ͯ:�Q�!7vn�\�����0�<p�Ĥ�16�6��wZ(�w���������n�,m՞H���!���-���x�={̧����Fu��M�����]�,N���E��F����T��]��U$�v^��i��9+��~�� �&l��A˥�rU��� |�����G��s�dGɬE���wָ/D'.�::���,2%��&�G����#���˾ȇ���o��M��e�E�o��<~9xšj�@�p���}-��꧅���]�Yn'F �U�JyY<0-s�����`v�\�D�����3s�g�S���m.�z�i������:�-��8WI���ݖ)a95�+J��Xj;�R��OkY�I���	�֤�kh/�G�>	��T�rZ��q^���Jo���I/�W�G����s�K�Shd�m��9÷o��=a�/�Z8�(���{��#�����Tg�3�m�Ȥ�r��Nd�Q��K%V�x:e[0ʑ����a"�laO,W�IǴ{8?�%ݻx�]s��6"	#���IE����v����Ak\[ey��F��x��e���ޱOV[��_���k�����=�����v�މ�^���Ҭ ,���`��+
'{���-ޞ�߃�������r60��ݠ��l���tS?�Pq4��nh�O-.��yS^8�B��7���	^}���}v�H�D��e���Y����p�I����I��w��������E�̕�=HRd���@�fվ��Ju���rd\�yˣ��b���L��û�<�I>no�sVB���s��k������&Q�Jw�
�E��?�\����ε'���D�l5���}џT�mI.k�T-Y�٣�s;� �:�^�Ö��R�^_��n��<�n��������3Qf�������E:�v�o��Ȗ�,���`�r�v���|<���t�j��t��������۝�i@Ľ�w�0$��Ht2�D�18�D�z�z_ ��N�J��\��H��"�7���_"�:�%���K���)�D4;J�1�c��#e��ί*�LM�\���I�׳�<����<٫�a}��<�+Wv<�5�5KJ�����O(�#��y���� ,t~���y�f�d6f�AH{��G����i|�v��u���x��F(4/´���r�Ĩ���哧�^�͘]
�?չ�B!�n=��:)���!�^��K�3��=�>5����p>N���H��<<�����q�?6�շ7i�#L0魮�0J=Hc0��E���B������j��>�o���B�G�83���:�);X ���3n1n��Y�@�!�pO�}�c���ǔ��yu��'�z�V�������e2��U����WU��G�bМ)2O�^� .���_�2J���gQ��Q�wX�Gj|�5�����]���|���x��' ��!8�
�����t��Ý��Y�"�a�7	K�&e"�E��-�ړM���|<��<�k�Sx��rj枓�v�Q��Ysj�G�t��{L}�S�3k��2C��"^��S�t%QP�˟<�Ifr���]���]j�ʁ���ם��_�c�1I���5YCA��A�N[iZ�)�a��w�BA���.p��L�c�(���?�5a�>c+D�J�&�Q!�xQ�I���b����8���l�w�:�S;���3���(�b!���s��k�u�>3ƭ?P]�6U�1ZU��`@�[�"6.ex�����^���NR��jm
�t���$:u����9�=�l�����7����Xy2��S�n0F��x�`�ƣO�hR�C�h��;S^�zSc�Hh�i2�`�|��M�"���揼���gCy�/����8J�'G������g�ܰ��)$%����&@թ#G�f9���栈gf��Z�S�	�*Hw]����[bU�z���1�W<`n���#��2��c={��D$�����|Z�F��H�̾�ܑj�k�sڪ&��Y����K	B1p(��'ϣ����=��~e܀l�}� �*���mL&�ɲ<X��r�Z�z	�%!���K0�G3����Hec_�^�q�b�1��H�!��`U��+����B�T	��}���Zqp��\`�~Sͬ�Ԁ(Q-fd���ڡ�Y�����Y�b�	�����b�X��>�L:����j~߶ӜS���|f�@>Α5"a�x�/�}�<�
�31L��Pp)�����xTq��9��4� a�@g�E�҉S?O;أQL�y�|Wt�1 � ��ĈQ}	_����������� >��x���$�oL~����i㿽���Nٛ��7���u����@���Z�Zs rj:�c0�D�|#��� ��D���&�<�?����l�\�A<���
�����y����L�4��b���K6͵p����];A����&��A�K��ꜫ��'�6��p~R��9�炸�22�B����9��=��n �z���ܹ��J._^��>�]S��?�M(�A�T�fY�ݹ\�/U��-���ђSg$�ٲ��k/�����iũ;�`�P�ԕ�B��Hc� ��X���N�F^�u��;�a��9���&���R^z����:���LD\���x��{�5�]{j���Y]��"����d��.o�x�]��*���Џp�Pc_���<�Cºp�ޯJԳkI{� ��ԥ~M�Y�W���Qӑ�	8|���C�)�c���(?M��C�i�x���R~�{�pf��8t�F5QK���!\2V��ڨ�_x�<Ǿr�CZ暓��b��7�Oa$s���������Ç�u�X�gJg	�;L�yL�}�c��k�a������i�+�c���{�+�ڃ���s�đ 6pg""��i�N�׼7�S:���g;�x0�R����
�޿�Q"|�6�ո�"�t㠓 ��4�RʹZ9,U����ýB�x�BQ0�RX�l^���]y���WQ�����o6	��"km���1���U,˕ז�(l��.5�G�Ə�1B8��ӮY3�V���v	����>�m���F���	��o�v�H4~h��lLb:���S����@����%v_�e{�{0J�pt}o(O�J�,I����b��_6�C����k��8�
�V1ɼe�%Eս�3 �hp8��̊�f��!��	�\�Oc��#�Ƌ��$e�=�������}7�I{Wl���Î���+ oVO�������W�k��A�.�{��������J=O��kR�f~ޓ��H�[��W6Oo=+��j(�Vc����pr\k��B� �IĮ��;�U�D�R�I����Q��(t^,��j2���������ܕ,�<�uLaN�O�c�>����?��wTF/#�*
Vt�z7I&��)���������L8��Y��J�WS����&�I]�P�3VS�n��𥩋�{j��p5�Ke�2�F��Hw�
�Kx�|Fa�ٛU�tGn}�#z�"$�{���֓7lǲ1n]�2(�H!�z��7�΃Ol�g Ⱦ��.� ��t�}�r{A4p�Nn��1�=�������ndkB Ѥ����
G�W���QO�\L�>v���G�c�جmA���m�D�kJ[�S��p��p����Kc��f�[	�5�x��?A��!�ͺ����2�[��P�-��C{\���6/��վg*h��3@��kUʎ�N]����S�'a���REu�P����v
L�xi�ݎ�+O��y��]u�K�n5ݺE��yy�I��g>�N&�].��ڦ/^�g�]\��,����GXQ��ɗV�Ȼ�{S�~J�dx~�d�u^-0d��snB�q6�����4����S��i!��jv��	oN �d��~X�vE��s�+�w� x���U�r�̆���oFN�ur�r��:��x��kN�m蛩#紐��v�O����x�����G� ����
�(al��#rV,�YU�Ȍ��ﵑe%�R9����+���kaʵn?�n�!HQ�J�Ӏ˫�����\�ո��l��&L8��o��/�V�_$5�V꩏Z4�}+(8m�i
���*��(i�}S�`eC~���1Y�SrbU��Ęt�M��c�Zq���:�C8^�W�^^v4|��@:��h����	��"B��N����
sZ�<���U�~�Ҽ0��sYc�OoT܁u>�L�~�rWS(G�>�Å%=�_���z~�����9mw�;[:�ҩ<�� 8w�#�b������7���4��ݙ{����%p��\�%>��}�W*��B�咽ar�uog7��|�2E���m�`#g�ށ�N �ر�f��O�1P��(O�[��|��=��i��`��9�ܞoi�ER��\��bIر�9�j�B���D���"hB�W ��DӀ�����!t��s�p�uc� @��(�쌉E�J�DB&���"0�ov���H�rө�m��a��V�ϑ!�־ OE_�̜����B-���N�x\s�&�K]Y^D[��/&G)M�~�OSrk�א?3��Ԣ�?�^�����L2�;W���P\�P}��{����|Z���*k�����]���z�^Ew7ܕ�e��}�e|�q��s�,<(��/�w��E3=/:�T+�Z�&A����ϒ0��FA </��Z�9�FG�������S��H\����
Au�F=�fԊ=�Ě�sy���@#H�.~���D�X�8�4R��x�z<x� ��^I�$o���#^Vƨ��l��<E����X@������L�d������M���|õ�<�ms���/���g$|�鿺������ef��u1��N������\�8�f|��8��1{����v�H��c�g���˺<�ʊ8㟯x���W"��ʜ˶x����4.H?Q/;:�v,��β0�,����l�te�9lU��>lZgⶲRg,��NI����O�}��z?yƋ���!��ꘟ{��yʄ��x��#(���Ppiʄ��q s�A0|x�nX~hN�����֬�N�>~�'ы��5�˃1U��EW���[��fe�MFF�yR�ł����4d���)�=}d�*_�ޢT:��oGvɀm����)��"�(@�[��D x~s;~a]�vm�ɚ(�}��||��G`���j
��D�*ĉ���pΦG���0�LNg�K����;جp�ˌ�=iob4����z��Ev44=G����m�ێ���_Βr������� ��N���p�#�r~��u�6F&��Y3�y|[5�8����{��u�����Xr�h=�V2$1�(����ܑ��8Wg"�XLu�!��6��u��Y�.\y�dG�O!�ҥ����ةF���1[�d*$x�V[A�@ ���	nz��v���{�.ʝ�pD�����^�u}/��0��G��@��<�ʡ��Z[�c';�ߚ�Mxrt��������Axvb���D#�S���41a3�ɰ���P���:Q���r�,B��u0�9q��c��bm�Oh�뚗�^�.rN߮2�-o����V��^&ƚ	�N�k�A��UґP5\w��N���}�w@W�O�#�9z��]�٠>�1��Qw�,���/#����M������0��q;_@���E�|rH���c��#�X�	9�Xы!�C:�.M7�TqhS���9�H�ǿ��E�����6U����({:��_Nl!@�!����>��TĎ�ɷc�t�W1�B�#�B�Z�'��t�|F�֦�E/[�����R���"�.R�`ii���R-��`����&�G��`�7o֌�$n��3�*cc�E��Z ��BkG܋p��b㪂�`�4 @p�M Xpw$��ww������,����,�����M�T}�=3�5�4�5��nړ)���6��y�z�������v��(oDY�7�����>�]��ʜa(n>y~�k�'�Yd����f�J*��D�Z}��gI�,�K`꫃���A���F!v��@2G]6z6�R�̗��]��ýl����Z���\b�Ot��!���^v�>pt�=0�NYm6����}����\i�z�yҨ�W�_���'.0�C��	j{���K�`u�m�p��EF.�,z��ި�(�8) �;���Co��U��I�V@����o�Vj~�����k�R�M~}Ĥ�2�Ⱦ.�a%�g�j�xK�rv�y9��.���Xx&�?�� �'Vb��I�7�!�e*$�+�߀���5���D ��0��)|�^쇲�xU*�0a�d���Em���X��!���F��ޑ5��!ڽ��n�R����Eݿ�}��y��\sEՍ+qZ�q�wk�}�!���A�����Z�k\sv���_ec%���~W����F�v�v�ݟ�R �sf�Q�-4`Weh�W�s�X=���t���X��А��Q8\4����Ǔ�ݸ҂s���J��|�R!g��A�|�L���Z����ӽz>o��j��%E�f�бg�<�<�?��Ģ��΁*�8c��YI/�vna���r��Qd�h!LlM��Rb�u��������ɿtq��I��ﺹ���r��4�E{��#����ʹ/�	+q���Tm��f�6?#� c����cb_ݲ%�glu�q�JyK����E��O[����)9�VZ
M��'�KtV����fx1�S:OCl�K����cxH��cWI�]5��@���"G�%�S�K�����M�&�\���%Y��xD���Dً�$<@��H��C2�S�C��qoq8�c�(m�삞�L >��O4����;�]fm"+�a�)"z�\v�u�K0ݻ7�H�X]Rfo#f����$u[�_m[Yg=�NrEmi��^��H�	近�"���Dו?���3l,�7ޗ�!�-��Kr+O�~B�����5W�cdՍ[���:���E!|�'b�:^���>s~���O��J��H�Z�)| ��f��(���j�Jw�3���ED�G��e_߁���Q�,��Y��fRYJ2z��H���!o�eۢ7�0T�`ރG�S�u1|;�a)��7�K�3��YDe�CΊ��7�V����yW�f��E�yo��9� �v����v��=Sɼ������i���Q%!.ƜSU�ۻ����S*-������͛{�>ش�����8��ï���Y�����Мa�a���[@��k�u@�B��)5%���rG���a)c��by�e�]EE�f��U2��(��}�^�Ɋɲ���8����WC`���)֙�>����L�6�u��5\�ȶ]qZ+n��Y-���I�n�Lz��|=KoN%\��E�ጰ��W�J��X����z�刑4o��oLRn��~Q)Mv�Lk���SX�U������y�%|�K�� dY_5�x,�ژ�i�x<-?2����[g��b���0�8�ު�{�\M�l큽!���uPm�x�켻��Y���=��ץ7;EZ.��	K����[-Ge���@*��:+���UY����N��(�f^N_=�w��C���J�w��҇�Zy�IM!~�xu��\�[a���(��čZZ�93���=��Ē���:�H$����T0Fl���h�.;����Xw4�h�k�����c��6���qj�߱``S��@-��z�@_��m�����Ty����^灯C�
vZ�!ϵ��S,����_�Mֲ���whHC �xV�(|�ߥ����*56ʉº~��@�w�k�y��r:p���A��y���b<=�G{ڱ���f9��_����t+-h�!��ت��w]s�����D��m�k��S!i� ��8�ҩe��Tæ����u/��P�N�;敗���^�OyQ<�D�4��o��=ct��[����2�O�bR�}Im�q�A:��a�؏N~��C.�%����o]T��]�fq�-�}�F���'9��`:o�<�!5�_����딄IX�(�g�:�&$_�"�-��?0!����=G�j��eL�^$���Pb��O�f�X��Pi�fL�LQ�Z~h�w8�L�AZ�"�����_�q�Ӿ�tAL%���*x�K5|���_n����Zo�큹���"�;Z�`o>Iȓ�������6����S���n�l:���=���|������8{-߾�*RN�T�����*��P�����W�h�,ci��rM�l^�Os��c�Dx��0�? �����ӵg����l�%��t0䎔t��������½�^���Ny���S�K�E-�C��+m�̶�^;.�&~u�+�6�t`�e�Q�B��r�q;�a�fL�m)�!��ܴ��騳5�"��������N���0/EZPv����� v7��`&������0�R���dm�����������q��,BM<�f��&x�f�q-;�H���H�8^tω�^tEà���e�+�ǾX�B�����N�J� �:����Õ�z � ���J@��:��wmP
L���\O<��4��1��w���<;�b��;����ͽ�dO~�� '�0,G�T�c(��2 �(�6�!C��'�ѝN�10�}hug6��r��/����ͭ�ϲ���u]!��I��V�+\���p�.1�mK
��w�ףy}���3�o7^�-r�����[�O�)�۸4;�8ގ�b��1��0ޖ�n�u署��q����g�/�*�]�[1��	�@�?4	_i�G{B��C�d�;�+0����3��N?��1��Y�����x�K��RW��0~�o�7�����<̯F��q���A�+q8q�#d��������:Q5o4I�'��'�0�.��-�bQ'���g�6��-J�ч#�@0�JX�gH0OVFV�����˟%P����*���_~b��b�|��s|U�o�sc����}q��z��,��V����Iv7���O��@י"���J��T��$��US<nkn삳�?v5f�O�g~Ȗo�$Ku8�wP��Z/�2�³_T�a0b��L�4��a��÷�t%��')>{��M9�sy�T�����Ar9D�x'y�j��L��Gz�u9F����7�	��?��a�o��D���=�[��Df�`3�Й�l�9�������f��2dD�g8�=���1r��،WlH��v�S1	�f]N�M'a l�P<Rƈ�+����ڋ�|>q�Z���G����尬?]���j�׷q���j�\��<4��1���ƞ�;x�H�V�tY�*�����A�
�t��0�jپw=3Z��n�����Ϣv6������d�@�##�q���xư��`r�P2c�S���3�BDI��O7%7&R(Mx5t�M��U]z���o6o.��X���v�@�׍��5�+�(�(�An���D^]O(T��[Ae�k1;�+pTT�����V���3c���a�Z{�ǁ�����Ac J�~�Á;�}���W�wa�o�ѫD�PѬc�k!���[���+��Ӟ��Y-)�_�O	T�4��%􆳞�tͰNU����6�՞��>�A�=�F��YZx��ʇ��9_�f�+�<A@NI�9�����OGg�[�����þz��lڃ���L��+6՝;�㴼�p��wS�zx:�f$�V.;��/ �O(�H�Տ.v��.��}��\J�#�Ů���wb��?�� �>,�()�w)��/\*_���a�,:�Ƶ<J�A���� ��[ϖt� ����O��dx�v�8��&z���T�ձ��G�����z�E�?������t�{��ũo��4�����m��7n�yB:-w�J��WY4F�$M�=xz�	{��*GuNa��c�z�_R�>��ye2��R#��O��wϖ?1�8\y娬�u�4)�+Ox��M��}ϋ({M���?bf�>6w7����H�x����n;5�������Ǧ�P�9��Ě�^��S�`+�=��F�}�S����m2Z�G�x����f���&�����w,s����]�Ik��)p�$l|?f�.rGq�����;�qɮO&b0�C��d�[��ؤ3��g��/�q�:�����g�E��Հ;�m�u�ɍ��ׇ�>G�{����ۖ'���џt�>�7��K�f��jn�q3���_љԥ����t/0zͺp"��v���(r� �6�&���O�"��7�WJ���?eo��p�#�ƋDP����u;@�|���f���N^w
�FN7m#�sČ�)�]]'��͋�� �~��sVk���k�>XFx����.�hEo�v��w�q�`��pg"׻�iK�w�O�����H�Y��/ʹ����׌N{W�6��w����:��[@/��.�O�@���36�/v�\�b�uO�y�?g>_����av���Gd4��V_��Ցh�hB��l~|I&\I�.I �`9t����i7S<�[R�����7X��Q�O�z�6��ȅe�LH3Ǡowd�<-H�h
��|��<�s��U��#g��g!ǋ�`�f�FTΐ�ui��Y�f��0q$zk*Id�xW�2�#�Zn1�P*~�<�)j$y�P��)J�1�x������Ȃ���d���j��΄�r��[������~���Q��ph��k�/�к/\�'QK���M�2}�Լ�Pt��?Y8Ob]�_���S�\�`��g�.�M�I�y$h�+c4d�\~�ͼ��^��Xf��^)���B�P�ny�$��JְάǳQ|�`pf�䫐Bcɺ��qNSf�q�H��e��8�b24�c�(\l�t�`�s��+ϴ��`���`̕�܏h��J�J��������/�G�[�#ؗ�bE��3���e�J�r,JRkP��c��F�y���+j���\@4��_^E�\�y��
?5����1LI[f��K�ǝ9ty��&�MIņ��DEzP�ej��j�l��p�î�W��$��s�TS2qҳ��1o��&DGj_��h�[�������'�����)d�s"��|�'��Q8y���4/��\���֙��>7�FB�:^��1�U}�Q_͜1��#N�����g{k���?�� %[����[�"�Nե�����-L�	ދ���O+j-�?�q�a����]��ʰ��i'�����,E�?1e\�HNؽ������Co	\��ݏ�r�ʰ����g�fdp��E�"����Z� �
D��U�?��Z�/����/:�:~�������D+�SpV_���1�vh���-��z�;�?/� <-r�_�4g2X��},`�_��#�����!aз�u{w���qw�5��`q@z+��_�(	o���1.�ٰߍuۛ�bB�12d;t]�B}Q4�tG���:O� E��d�~�}�]����o��b�m��j�������\O����_���>~T�f�E��ϿΦz�Ƴ��4��[��%�����r\�8�F��m������=_9�]����}��b؈���A��q4CY�1���>�,<�?��/�+h���F���C=��ܡ�8xO��4��~{H�+���]Zzb��u�+����\�{S�\�<���u����2`�-�aOkZ�{&���E�Յ�e��Dn_����Ź4\��y+�L��Э�,m:Q5y7��4��"�#�ţ⨣�+l4٤l�h좕1�ѷ�>�[�i�r,J�ϐ�q#�q�?�N�N
9#�9eð$�PyZ�V���XB`Sg�{D?{��R�'M\q����j�R�������fT=��ٝE6��_傶�Y؋턿����UB��&�I����Pg[D�0$&���H0t�N���k��PJ�Vj9!��+�q(-bQJo&��`L���-�����9Iq.��6�#���5����j-���)icea��*��=*L�*t�H��U>�u���J��9���2E�l	�l�
�Q/_k�S}�d�e8����Dw7	Hg	�W��8o�����Ng`-d�L8W>��\H��V�i�Te轗J�D�q��aw���+&���}�Y��y�^�K�,.�m������B�^�X ���|ٔ.�B�	��DI ��7�C`����8U���k]ߎ�lX��K,�I�YI�~���)�N�g���j�*�{��K�� �� �cWm��U��Ꙕv��eJǹu`��̪�B��}�V�-vۦ;DS�}  ĩzZ?�!�����ߐxҩ��ӹ�oOZk&t�����,����������%��1Pn<z��H�/z}F5v��8!����W�eh�ʙ$�c����ݬ:=�L�lX9H�|i���Y.:��b5�T���4���������	}H�Dܷ�K���9w���D�!�Sû_��f����׀Se���̪��W�F��1~/���)�gq��N�8^�m8��8�������� H��=���i�:�@t0���>T�
ipml��O�6B�P���Q���R��P��/A�x�a�Є�����x4@�X�!��Ï�>��@k-�;H�5U���_�W�a!N�r��yD.�Iei1�hQ�ڪ��ɱ��D찑����}p�J V�c� _b ;�/�ÍAd���>�����)���F�O\Ǻ�p��ѰJ��p����J�Z�yc���@u���Z�)�f`0:�E��h0���e~(��:�,%j.��8%;�Q ��$mlǴݙv��X\O*a�a��������
����=|]	�BW������Q�w�E��;��}/&������&M06S����ݯ���X���#-����L�E�|����b���Z�-iU��vn�D��J�~��>i��T��>���J���/j�/��u����w�F҄���q����������颌��q��E]7h�۩4��WrI�S�u6!T�۳��5�h����oul����	�g�8}�8t����4����5?�e&�&2�Y�9r��+ʴԟ����������5@�磗-xA�KtS�Ods�ۣ���ͩ�ەo�{pb��{UV[��{�f^�ε�֫�,�:����l���p웉o#k~�}W��.��>P�EQ���������^x �兣���P�-q@Hq�0?'#}�R�� �y�>:^W��?,��C+�M:��M��G�0p�z���8��U*Rp��>�J��w�$+ra���;���#E�?F�J?�9svޏK/f�"���Fb�6�����Z�/�K#��s�Ͽ��4���� �L-N���j�ITQ�r��~OW�Ɏ��X;�����Z�C|V~�r�V��+�G���;r�G�&��(��������0��|ƍ�W��~fY�F�fd���+z.��$�_]���4�Ǒz�(/ U\���p�~���Dj��=�ן+�ph��O}]�W`V���#ݼ�v�<���s�T�'�b�Jjy\�'GN�A��&�T��	�b���F�ӊ�R�hj���KPj����,�}=2%7R���4$��iI�'��ݏ�
�Sy�~��'B��k���m�|����F�T��u��U��	�b�������%Q��T��3Bx{��]�)�w�����M���w'?�ς�2��Oj�`G|�/(���V���3���$]���:y6Pp{�:F��.�W0?v��x�vEBu��;�\��j�Ҿ�m�LV���<��5�_�-c�����xه9�e*Y\yۓ�I�a���;
��K~"�>L��-��6nD�m8�i�������d�bA���Ѹ�p<!Q��y5��vvعw���!ݛ+��%�`ՙ