S�|��8����
�>Vi��-�ba`g5�a�]���6����(i��ԍ�2C�G�픇r�	������d険�R9�z��Q�Ѥž�*��X
�'�+�*5�x���JG�����dT9I���W���.�ÒQ�hz�ƨV�zI�[�.A�������o!4�ᢾ��'��W����<na\D������G��/_$��n.�q��$6�dB �X�����'9��l5\�]�,D�)%Vm����T���������)}T���W,-�r�\�C,����ip��c[�5��i���.�R�+uH<���x��4]��M��x���E�`��`�Q��hEm��tGD����d�����'c[�ʿ�2
}����ŔԿ�R���Φ�%S8�G��^a�����P!�������\�~�G�~,�q��(�ŉ!���۸�qU^������츘J__ ������B�1��܎���;����"���|T�ј��}����4�����n�޶��D�K\�`T�H��7����5��n��@����<u�9V���6O= l�p��%5� nYO$K��m2_� '� �]�h�`k��ˬ*`Nd$~ΰ	W#��K�a���܍��a��٠M͌8P��N�aeY�v���RPW��$#'��r"&e�1)D%��G��Mj�C^!�x�`��)P=QyO����k��NJb7����)�bJ��n�E�k]d�p7
׺Ѝg��1c��Y�H�۠z{��i�24OK`�7[,��F#g����9��m�U��������Q8B3=�(��F��+�U��nu�����z�[G�a�i�v���>�b�fw�����E�Ӽ'Mx�S��i�1ժ�y}���_� N�ۈb�庌h�d�/n�L�+ک��S,+�U
{�F���w�4���/�'b�,��,��>8���p�n���:y7��{c�C4U5�|I��vG#5�(�-�ܝ▆�'
�����` H6���kOChk*�Q�����,ԑLGQz~Q�oV|�����l��3&QVmf�V6I�eP�za8����q���p�<�4:R��@���!A\��WF��8,@D-�W6�^}5˓|瑘zi3;=.��Bk�� ��P,� �W�A�r��u8r��ѣ<lV�j([QV.�
/� ~�������p��.��DAA~Q&�˰��5����͕��b Ym`Q���ӀE{47!�.�yf��I�qO�n��EF9��Kݶ���$�G<��Cȳ�]r�Bcn���:�>@�)��}#�� 5��[`�q�"�`*:�j2,1ޏT��pj��r�����&�#�	e3��ϥ=߄ǍȐ��k#G�AF�ıy�����F�g���WI�?ޝ��s2нQ��5��W&6�1�` 7�����zA+��x��y&��!��%T���1;�F�K�,M�O���	*��"�#u��V�^�|)�D�����d��{���� ��x�[i=�p�`�*���U(
��ν��Wg��[Ƹ���U�s�_1"@lWK��0I�