q���{l����U<	�����>^t�G�F^<8�^�$2����&1�WVn!W2�"�����gpRp��EW�|E$%��h��Ա�.w���+Hh�v�9��q�f�3:i��]�\���:��W�����a
��r�
�>�/����i�3F/��m���J)���󜊡!ꮾ�v�u���	��ȷ�b��ٲ(K˻�/�F�-Ռ�'
y]w�G/��B�	akBh=d=�i*qi���Vh�8qnɗ�K���E�1C?@R"|*�<�^|m
�9xQ�m���ADZ9�v�k�cS�2.6�Ʒ"�SOk��:�=�D�d��PC����#`�t�sxS����2�w�Q�)�;'l���ߐvy>j�s����o]�Ϡj����S���'�a �j2�dܶ�����Ti����wxo�����0|L]O�^$-�ΒV�I�.x�~��Ӆ��PU��J��� ϵ�`�}��s�ÊN	U~��4<��|k�Y�!�-�R�a�>e�C"�r����r�E�O�.h���n/;ЧS�����^hYܒE!��,�h=�����M�G��=h�K��?��-S7
�'N�� 2bl��>����&�$�I����C���Q�	p��ҒB�'y�.=�^�v !�,�k��єЊ���W���~dL�I�%%��ٽ��	(U��Օx�����U�#ub�E����u�S{,z��.�bw��{�R�rr�Ƽ4��o�/���`���ǬZF���$Gؚ�7�N��Mܿ�,}��u�0�k��u�0��ϻ��5j��_B��Y�;BS�5�cX��ZQv�[װ���4�d J��Ǐ��R� ?�6��U�3���e>ˬmO��-��ڗz�T�2����u�,n*vo�##rb��`j;�T�i������8A,jy���h���`(m�����}���@v�E��<@)df�����K���^ t�
�"�R����S�W\w�o��a�4�?�֠oErͧ�(�&�Degv?�q~JS|��
Z��zM�LJ˚"�`e�d~��s
�9�߾{[��תII�,\[֊|]�+��=\�,#�9������l�ʱ���#,���o����@�Pq�S%��u�����srLZ��ۆ䆈ad��?����?��=��Jh�Y)�"_�Jh!�����HJ�Yl/C=�b����Kҵ��D�0���>�������O�e��;U��C> �"�S_My�sl�܌���7�(���˘wg�'��}�g�Ꮓ�h��,ą�a6�m�-7U�~���r^�Ӓ)����d`<~���!����f<����ߐ��F�І���Y��������*S�5e-槨���Ą��+�C:���(V�P��]��5��u���_�`�݂Օ���[��g�n�-%@񁙴��Z�}[���dG�bv�*h��؛>��w�ă8�_�9��j�ȥ��=��Pz�v� tKΑ�4���m��l���.�E�=z����zװ�N��}��7�L�E;�=����ĝ���qIJ�$��Ε��؜�c������������5>q;�я���[�R?��(��V	%.�Q��@���ĳ{ULҍD�-�ե(�&��7��d� 8��i�����w��VO������=�l�ȉ2��x��c��N{������~����e��3Nx�t��?�j�Zm���t����H�P���"P��׻}7��SNMق(G�x�*��,1g��L����6��Ex�x�+o���}��P&F���j��F�����]�,	�264�~�L$���}Sw����J@������l�w�����{�qj�D̩�i��[$��.�^��1�-**�����r�gh�f`3ܜ��2^|��"�zM[��Ь*�(���։ñ��>S�x�{��m�#�U�^w�D�{J��_�Y`�q㦡�|�hRNC��Q�3SO��)�2{[�7���&�K�DGJ�ϖJ�`��R�[�qg�R����:g�v��>�
�O�^�ߟ|l�%�Y'p;ݸ���N��������lrmmc��vpz�uR$ ��iL+p�5��S�V�hw�B����8
�/�^*:w��F|�c�~L�[w�<0����[�M�Lߚ_l8�O���
9�՚S�/'�q���f����K���"���:���#�p����?�n�����	}��^�7iR�j��=0!\��7��$�35[b��l��%��z��<_��l���E�*M_D����ƢSe����W��=��7R�^g��](c��,�G�e	eh���.H'�q���_�չ�z�K�H�zi�|����qLynL�ni�o�������>U������3�m�aܩ�|���`��:yS7~���<�)�6���DL�mSCl�8b�M�9�4;jbwA=e��|A�ϥ��4�&o�j�+Z<�?�W�]�|�����}V sJ�(�nӇ*@���V��8�w��H��am�Q�?ʌt��z��C�?2!��XL�N3i�}K���͘�N��2NK�(qO)Qt��0��?���ǽ�ֽS�����H�*��v��Ջ�ԽOM�b�i"�Y~����.�yU�Ħ�f�z|��������ȧ����x�+�麬kQn:q2��n!Th���;E-���#�b���t�؛՞8*�]��M�8�Y[�KK��p����2�[��f��bM2��mC�q5�[Pȁ`~FgG�Z��?���55�� ��+�=���e�`��œ����p:x��f][���-P�z���K����r�/+��e���,gԝ��M���n�}��.�P1u˴fz�r�1pi͈��b�mA��
�-j��1y��,��I3Fn�w�&PШD�JԾ�2Z~0��+����L�����l��S��P������U�y�ҽ�8rKc"�zZ�~D&��cZx#2������1'�=�b�����h�� ��[�7wDs=��+�ũ��gm��b�on]�/	��j2}�{��]�?MPp��}Hs��ѹ����C�0�|8�6j��Ra�D(:4�;-;���+�[o���@d؇a���m0�������Hk�?�aI��WjŔ6k�|�����t��y�L�$;-9+c��WǏ`7�쪥]��������+$mbW�RkIO9mNԐ�S�^��k�_�Pg|���C-ɶ����ޅ���F�{&ɯc�F�ޯ������q�8��>��#�H,��Cb8!}�i^���Y^�*���^�O���LSe.@-Q�a���RN��L(�q��/��R7�|F@Hv�z��ė��W�/0�f�iH��6�(b,n�[���Ac��ş�O�����U��bc�^���f�W�)�&
���?x��!���!�7K��=���ּ� T��d�>4@�8��z7��^4y�ݏ�l���=;�?l�� ��I�4�R��Ͻ�I����NGf����߿���P�Ã��+�|s��]��\�P������uŏ�,����)��M��[lC3t�$&���Kk�U���{B�D�4������0'�MYХ��T����P��=�(^΍
���WB��I��#�?�����v'�