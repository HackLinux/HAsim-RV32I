�)��o4t��a�z�&��'u
C�a��۷�7"l����!'�?+i��>0c[��6j��|�m= �	ڿ����ho�>���T�d+��|��Lď+�Y�>�Rh�m|^5#u�#~��A7�	��Df�7��&���!0ۤo n�1?��D'|�����-p���O����U�A���&��[�ے*�=0�3����rb ��Л��z�������,8�{5��dQ_OGkb�c���d�cɚ�[&�jJ>��n�-#c�`?�j�!�h3%p8K�<� [�nئ8ZX>�����		�����&�YcR1JF���D��0nD�+ N9|������<�8;�&4$��Vw�&E`��$����B�;t�>E������v���� 
�ʻ�%�H���A��UC*�(�a^%��a6�[=u�2(2��ep��y�9�)���'�(߬���/��P�+dZWV@y�b����ƭX~5-�[�Ӂ��,�yRh���ǢI�6�q�+�P:�iG���lF�����l�ZC����.�m�u{6B�j�����.��r�Y�W��WO�7G��!��ոl�������dC"e�}T��)p*�oȠ�n����܏'��S����q��d���9�{zi�:\�d��
��j��2������T���R�*�0�_�i�D���/r5�d�L�&xNa����UX=X���eË�Q�Z��᭤Wi�	�|�1��)��C�,�f���UQ;�{^y3脶�������t�O�,քHu��5�_>������HfQx2x�.MO��w-;����)���!+<9���&�K܊Q�`��
6�m#�~s�)�F��Í�����2�?��a���:7-�F`6k7/x����W�ɢ �@R�����&�i���/D�m�pr3�E�W�)4�\ꄂJ�����8�$��p(޾�"\�P�'럳Mc��.ԮJN4�1�=���L�G�Pv�Ģk��ǆ�
D#�U��|��������7��V�q�1�p����֊�R�qɆrE?l|?EEiU��Cg ��D���s�7�����/��i{��!9&��m�C~��N���,��'Q�7N(��J1�>Dӑ��=�Yd�f鄜�l,����}&�������n�$�Y�a�=�U�K���'&�hC�x)�&����U茯��.�����&��Q}?��z�L�634YAkG���k\��S��r�D9��9�ɬ Mʵ�����
��]�|7�HZ�|1(��M8rӁ��a��'�w�^�H)�������nO�_�Q�av�b5������gȯƂ��!!x�3�;7j{��y��V�U�"zd��d��n����s3��>��a��&@�Or�~Q���I�V�&�7���RU�� @�u�����3k��U�q^v��N_�2�K��v����F&ţ��/�'��󁅖^�Y$~����s=x̡�����'��p�G�.�+�L�͂����q�J%�U�)�Tu?|J\�*��/w�YZ5OR�|���"T�S߇]��|	����z�3�n��y�~m���a�۫Y!~G��A`�E���1q��l}F������N���[پ�4���L[���ww���#�,�\K3�f]]�Sg)��l��M������$R���2����U�A���5��L&���&�Ag߯pf���*�$p�8�n��;j�<����Q��I�h�^�[+�P��b�tP�����m�:�j:�G�N�@0�a�o�8?I�d�A *05I6s�������W��sڔy1��u~���)����#s�F��xgRr�d{��1�]֘O�
���o���OT�	��BF���]I�����`�����p�Y�!`�ހi&�!>�,y���%�o��Sm'�Z��������ꀁ~;��ǂ
�,����:�oګ�2��,�ű��:����k��$�bO�b�˽�^>��#��⡝^E\��v"o��ܜ����S�|�B'�15�\�qR�jz��)��A��|5G�
/�"���3���c;n��vfB��N���u�	�đ�H���wbwA�'°�(㝍�c��k>�"�rf�dIl[�(�E���A�m���B�w���"��a�w��!�TD	��[G� �"�y
�CK���tgV�\���GCd��!AY�+�~oZ.q��H�9s�F']�v�}a��}`���i�G�(�K�?^�����m=�&<����$����ڃ!{$��p՝��.	�`�K�s�\ij�j�uSiy�
NM���D=/�UGJf�'bv@2��$,~Z9��&f�*�,%c���f	�d���#z�n8�8S��� �$>�#�d�d� P����b�B�_�
�!�"���e�:�E�:Z�ST��U��CR>+�����rYP%C�gE7��~F��m��R�U4��@"����|]ι�P?�ڐ
qd���(��!��ĸ�)����,ӊ�Q�����;�A�������.n�F���@��ϛHC�x����]���2���%�d�!�S�R+�Oҝ�=���d_F���	��nc�|~���C5Zʖ��qݭ��c�9)��1&�\܈k���A��Qp�B!��|�i��� <sF��Ԍu��X�]�M>h�
Ǭm�i>�W�][hjѺ�, x