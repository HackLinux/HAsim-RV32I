5b2Y.O)E$="785'75)86/:80;:4>=5?@7@B:BF=DH?EIBCFGCEKCCPABVAEXAHWAIVCITCISCHTGIRHJRGLSGMPHNLHNJHLJGJKHLPHLRHOUISZJU\HS]GT^GV]GV]JW_KWfIViEVhBVfCWbFV]HXYJXVKVTKTSIROHQPIPRIQSLRZJOWKQTIPNLNKLMLLNHKOEKO@MQ=MT>MVFOVPOXXOYaMYeL\eL`dPbjQcrQetQdsQfrShrRhoShlShiRgeSfcSe`Pd]M`ZK\VKZTMUTMPSKMOIKJHKHJMFLMHLNMMTYMV\QXZRXWSXSUULRRDLLALH?KHCIKEGNDGOGGPKGQNFOPDOQBLPAIN>GK;DE7@@4>=4@:0>70>7/<6/<7.:6/;60<70=4-:0'7.%8)$8%!5$2$2#3"3"1"!0! 0/,, , .#,$)*()))('&'&'('&'('''' (!(!'(('(''&&'&&&%'&'&&&'&%&%''&%' ' (!("'"("(%($)%)%'%(%($)%*%+$.$+&*',',)*),(.)/*.'.+/./0122335554455475658787<7?7A8B9D:G;K<R=X<^;b:d8e5d4`1Y.P(F#<685&96*:7/<:1?<3@=4@B6BE9CG9CG<DG>DECCCHCBLBBPBDSEFSFGSGIRFHOF