���۔Х���vx��̝��8#��H~0l�bS�	IB:��bp�|�t{$iH	��� 0FI�I,д0R��R�)�����)���^�E���wvKC��{�� 7��8V�p�J�PUv$ A�BBcG�V��H	���m��Yb�Dw���m�[��)�����:P�g��_��r �`F5B��s]�V�v�l��J��``��~�$�\�X&�V D ��_x�SDz���w25�+�Ŏ��H��#�uV#��]���dݝQ�V_����$�з,e�T*�*��2��:+U��u���rX +	��q7��E��k��{.y���k�I�!�ܢ������W��n �Ȥ��b`����e\��   V��a�f��k7��4_i�x�,ec�����=��DԐ��0d;;�Rl%��WEQ���خɺ���N���/k�����N�r�+G��8v5Z�!IQ!%�hp@.P
�,�� $4W�%kF �V���*
�QX\}�i���bp��qz�$�\�"�pF -i�_f�%l����gY3,�>�e1�a���/{�D�_	�h	�|�]��=[�P�&�V/X5��h�� �BAkP;CV*Pz�У�hd؍�5��eV�8ې	t|��N�qW���x�PI���Ƨ���n��`p�
ةx�0fH@�   q�w�e�)$V�Q���U	��C��DNd��̫�\���������v���F���/h���\cV"11
������:�-���<d�E�d�j��
>�z��RƧ7I�ĿJ�z�JlC�QW�K�p��.���bp�usv�0�\P��0@��/��a[!4J� )UD!FqNc	df9���]�u�}ޟ������u����G'h6�z�X�c���frA������6?�S��	7'h�����>����"H-�p�܈��y����6ؔ��g�=�^J�2��.��bp�istz%"\��T0�q4�H57Y��0�$��s�摠2A��/J��?f�5?;S������`f� _�Q-��l�$(e�����52���RfNl�X�nF�&�����G��m%�&')�;�����Pn0�W��X2]	0���K��"YM��bp�
��tz$iH	���pn�h���_mS��b��HN;����Ŀ�JIlmȩ� �3��R�"R��KO�о��K���ǜL'0H�_�JF��W᥃�u=�3��*N�3F�ZV] Y6j���痨�������^�(/I�t�T��:��`p�
Էv�$iH
��� 0FI4�E��_I����ХH��VR���,,FꐪK�&�p��k�?��;rB��Zg���� 5��|��s��`eW���
+@�h�LMv�T ����?���K��k.��.���4eAA2�* ebc�(��.�,TH���bp���pj<�H
)R�p����4ms��sc��eh�������f����i�������Z\Xn�WM\���(D���X��Ћ��Э�D�*�d�� 4p��x�\_'��fPi�X���{P�o��տ&�V��IH�@^����7C^7�i�l��b`�Mx�%(\�`r�DHt�j* ��l�*�Qi��tu� �9�G<A*�TN�a:�=U.����zJ�`�����|�#e�0�ÊLlg��@���hs��O�D���@�����0d���|��ce�S.��&ԗvr/������:��g����bp���tz0�HHN�T0�(�\���-v⧠k��hqG��AE A��Ed�*�V/D�_~������֬����u�ҧ
`�Ј?v�y=�e"��Ľ����{:�B�M�YVj�q�-�s0�4�(�r���Ko5�fۑ6N�_n��3L>��-2J����`p��Ypj1�\!
�l@�q;�9��l[]M�ٚ��z��r�
]Z�7�F�=���ѽ?�)�Kd-F�2��X�������Ȭ
�SWw}���گ�Ѐ֫`�V��r�@�+J!�ֺ�j���uc,{�QJ�� ��I�A<"��d����ǃB�&��bp��r�<�H@��X(�q.Qa�=�*cL�j���tc�4�?��޵o�����)�Eٜ�f%E�_5� b�.�f�_7(d������_U��Wb�&	��Z�����PFoɰw-nKU=���b����w\#	�a������Zq]���~'��>���bp��st�1\�)�XHDp�v �}N$fv]�F"�V��V��Ȉ�n�������NU|��bD�0Z��J���b�?ՙ�Q�SN�G��UI+K��`������b[>�h�v�$]*e��f��\����_�5���)du�H�A����bp�-st�=%\�	�\0DpxQ���a��uGq�-.#j�%S���{��DuV�d����,8n�E~E�2B���7��D+����Y�`����%X��$�Y��z���Uk����F�m�5�^�Ʀsw�A	��Z�<�Բ3�	(e=	����``�
��v�<�H��(DpB��&�!a����jXH4>`$�d,v䋿�~�kr Z�r)6�,TuZc�o��/�ciIS�I����E\�8=g�;��[�$����vJ�k|O&f�ǶT��{�o�h˺A��o�5�;�"s_VOHD*.��bp�
̧t�0iH	�"� 8F�((��Ag���(y�-(�ˊ�q�/'�M�[�F[��Zx��hX�$�S����,\�4�M��|�
�Jm����#@I�W����}cB�ˤU���(eQ }޴��)�*�P �5���!&:�Em����bp�mcx�<�\��"�t0� ��Q���3f\퐿�ǯ^c���T�ov�^�������������,�Xj؀ej�އ(�\T`�U�1�G���Km�b����AN�aG��Ȼ���j#��Q'��j�6��d�JV���W�ʛ����#%���`p��|�0&J	 .� 0F�6��V�t����
֯ڵ�N�0�p;��E�ڧJ�4R�����������c*s�]x��������s=|��ٽn��]�s/]��
|������ �,�	�\�F���z��%��
�1�*�(�׉w�q
c����\����bp��up�`�\��.�XJD��pƲV�SnId��i-�����$du��Q@O�Y�VMg�,�mli������5S�P����on������s��>����˽��uJ�\�I
�C�q)k�Ww����Q0�e�z�����a?ə�k'�R�*I�1�