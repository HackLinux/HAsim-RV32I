�~�{��_d���M���4!�u����Ȋ.'՗v(tGT��֢I��4�Y��=~C'�ܴ��Y�{�
]<�oJ`��U��}�;�F��������̗����t�.��u$��Bd.�Wd�����M}����	(ϗ���BW�*�L
E�1�R\���?"[TS���FPP�� �/,n��7]��K#o� �s*�w�H�~���¾y���01�ק�����)�ơ����y�P�~t
��g����3(M�o5&��Jfgd�S�\�r�\կge�������y�!2e��	Z%�޺y�K�T��3m�*��-�E���(H��	��Jh�d�E�*���^{F��zfN	&��)12~w���{�[�Uz|+�� �OF���d�R!��ֵA,�x�d�)��:m��ݪ8�H]�im�D�|��kyPwzT9ů4!���F�	,X�0Sھw��0j{c[JW���xU���� �b�^fr�c6a�!(�e����d�wY�� F�v(a��C�n�����2b�W��N�H��7�ǽ�ל���m���ݴ�o���"t�҂AښX��K@�-U@��ܔ�����y�f������򊩠"���L�3-)�*j0����1����+��,����U��71���ԟn;v8�������0uv~r�|{^���Nkns�>�������+�j�
8wH�Ѩ=��-F��b�+u��ճN�s�*K[�)Sui���CFE4��W�;��v[._8�m]�d:CRJ��_��3Q�Z1բz=���$)�*y?�D"�5�N�%��w�z*L��A���ˋf�s��v�Q?�<oN�0�>u�3D�=���$�UaQXu�c����3��cq�à7�t~F����<�t����!�x�����MoV�ܐ�`�`�OE���M;��B�ar�Q｛k�C�m�v��N��NS���l��BC��S���mB�Z�8V�h�w��S粬���2u)ύkt�P�8����Y�;�
5��=�All+����s���g@m��h�炤!�z셸9��a�����ϙY"��T��҂@�[���qB���y7�H%�OV�cg�\�e]4��*!�AN�)�H.�2�@F�)(&��o6y.<)�M���a�و���"K���$���1�.�e���L�}�D���̉���@�
Z]�V�z������$��d���oJ����x=��MG�<��Jt��S�^�ȗ�����a��)�F��������U�P/wƍ6<c1߄�%".+ڠO���xQ��q�:d�!�TY��j��O�:p�ب�$3��߉�1����'Y�q�K��AǓp$F���GU5��u�ǧ�ߖH�����w�@Ý�@·�!R"5�V�W��&�ɍ�&D5��
��R 3Ƙ3��O2ZO�h�0ec�g��^vG�~�X�t	�R";1	}P~��lU~ٮ'p<@#Ɋ�����d��V(�8/�>�����.S���+���J��}�0�ʋ	V�H�45#�q�B~wa��w6�m�y�&UB�M/��� �U �=\�~P�����B�R����*M-�JzBP>#GK����mƧ\zl(�(qm�3��=�ߢ�s]�R��t���]m���)m��)@��JKE�ō�)�u���l�{a���E�F=�"�|Ѿ_�-���)�ȏ�+~�@��2d�ٶE/O8O{v���4MpN�~��Z�{�1ַ[&U�����7�P��4bKNP��0��ڑ_��q���.��c?c ߻,4��X)c$>䞥T��9�W�S�,rHߎ�V�ؕe�"���`$�Toߨ�+�/�7��hLJd'�|�?���m*H�I*bHG5��(;9k�����bZ%,�ӀV�pT؁3���ݞ![�%�v$ib�44��|w-�7��7��};7 �S�6=�)+gU�9ts0��wb/�{��w��WU�^	��CW��,��%���*k3O��Pf�J;`�\?~>�3;�8 �C�ѿ�Fo�&YX�żq>�|�
Y����Q���;���� �7���q���!�A���EN�HckN�b�긣İo���d�Z��h� <��S�6�V��d�Al�@�s�e2�)����D:k�:�g���p���\����f{��� �L�uX���ݞ��+�����Z=