ݴ�8�P�������k�䆳�������g�� ��􍢽�s`c�+\�=�{@%�)Hh�+�m���͏dI0��	B/X-H�65;��;P�{z����T���Lg�ۃ�;�/����~�����b^��bE��^��@Q�4y�{���nMMY���5YE
h7B◨L8݌��U��t�ש�f$��2��>:�vԔ���lF\�؝����X��˦A�k�83��xR�������j�'P@7 Z(�Ƴ�f��q��nZ����Z�^jЀ�#H����*�Sh2Gϩ*�4x\�f��v`x@=�l	��D����`@
0Z�L��'8l�?U����h�� ��" �8�A����O���r\���q%��XݴJC=�׀�Ci���u2�jw����a�1r�~�����:��Һ�;�s�n�Mdtb�xIus��h�wH�f%�Q��+Z�£��udo�0X�L4��{����N��I��
������ �����Ö�o�����r#�*[�^<����q��R�:�ѯ�d�0�n	k���u����䐪#�cW���T��b/�{��{`@1���o�R��Ӣ���RW]Cs�Jq_��i�E�?�rKK�դ���, e� �t�V��B���<�i���кD�6k�a��duS��U��?
�I�@�9�q���an]��҆�I����0���C%�rj���j
g$5T>��Y��0�ZjM�V�����c�T�R�l�������5�Mˍ�,�c	!CXqk��:�U|\l�W�#!�*s���?���IK��yGe����j͞��D��wN�����F�t�t�) 7�^']<ZH�lppO�� �c'�M,p��BK#����ɔV�L��˛jg���o���0eƅkO��nΎ�)a�P�W��j:�>��BAU�a�睈�`wB ��!� ?P�o"W��h��3J���l���Q~y{>�Ҁ	4��Vc��d&a~����H5u4,���V�M�� ����"u��r�C�BH��&0� ]"����X"�憐�1��{�P��m�3�.��o[��NI�ҔVV�ȀN�#�5��x )�Y�d2;�'�'4���tĄ8� kc������*�
�V	 D��D������Y�̜�.`�<�5��;��?])��9��|*5H!AP4 ��kQ���+*���e`�peueI�������J�P*-��Â�e��D�z�tW4��f��a�3�7�W���,W�z���8�9mcښօ��=��+"�)�0B�=(�UeM��U��xJ��x���������#e�I<��Afմ�M�����,,Y��t9Q�x�`5y����b�_0� �M�>��$_p�.� ��ȢĠ�!��y�<��wi�2-V���f��^B���:������l?�T�cT�䱆|��"���@.i�ɣ�I���çd��h��X(0�cr��j6u\Z�1l������}���[n��؄2��bE4H�2&�:��(5}�����,L�g1!]b$�7�`��塦s%"n�pZFB��E߇��Ĳ2Ama�V	S`ߴ:�oD]���}�cMM$��&�Oc�K.�Ai�8���<��60Q V�*R_'8Az�%��@���v{�?��sYO�?/�5o�%aM�T��_��Uf��������Uf�_���:�~�Zqc���6#�4 谌l-�R�oEH�zY~lE�5���I.H�	�[LU�ݖ4�gH�	�B��xJ�+/�~t�&��_w�����O0�y����\���d+�<uBc��bi���%&���)�$����Ӊ8�HA+�g�m��Y�L�w+YJ�*]����Y��R;�U�Ֆ�h���h��L<E�d{͍���<���s����u�v����I����#��a��2^�&q���e��"a��׃� �K;�`�����#7�6��g��\_9l˂#�t�FM� ~��3˽2>��qȅ���&���G�1>a����hYx�-WNjyD��'B~%e�'?�:6Se��.�C��g������}Y]VZ��TcaT��V z��xG�CJ%K��2Bދ�61��眞a:�C	�j��փ�bT��"�U���e���b���]��8tb�m��*ED���42� ]d�#z�d����2��j��]N��r�x�b��jZ_t4z_1D4Pl�*��ɿa���f��J4�����;��ˁv�-�� �`tu")��LC���+�k� �ʧ�W����?(�cSE�\v�qyA�3{WW�3S�<Ku�JA�%�;V��D�!9�$QH���:?9X� ڄeY�y=cw��k9�5��)ޛ��v佷�=D��ܭ]�o�kV(�P�����\�&P��
�=��Z��[H�+nB��t���jk2�8�[χ����6U�V?�a۳�/���&��+�������/���Y���ő�xLG �b�a��ا:C���\n1�����19�v�Q��5��ۉk%V㷇R:��- �#G�d�l�2����F�C8��d_�7%Z ��צ�N�s����<����=�{	�����I��	V_���N_����'q	v�CV����w��U""Hb�>��}�&7���1�_R�i��cbBI�2 �_Z�aA�i !#���� T�b۰P[�~�}êſ7^�X�6<Fk��7쀿��.L|�j����Y'�`��v崁�Nz0��%�z�3j҉eт���|�͒����7�ՕPϺ����^)�-�X细�j�ZM�$�����8��Q�-����6�k��ˍ�P�`���)�n�OL�ػڸ�pt�?�/����mr�]3���'�Z�����M����x�O�I�|���םq�i
KLP�BA{����{	��Z�²��r��X�}�o�ƃ�o)a�/�EJ
�`�g"�w���^!���(톮k�@�~�`�NM_v5ϲY���~y�	��ŷ��i�����fr_b�&��EO�H����2��ʰ�e�����`lzث���%̈��������+�Į��H���"*9����w[�.,����heH_���v�뚠c�i]�C�[ǜ<P��h��4J��(�.�t�\+�/�/%��ڒd�B,D�#�y��\��4oS�囵�4=�@��;��kݙs�j�tk�|� �/מb~���oD^L���=������SW;O�B{��*��t$������}�P?�����^�Q�����T���Da�����[1���^�1�[�5���a���w�$��G��ܰ��w ʘ��������i/�m��D/�R��[[�3z��O�����#��a�cY��2�ڙl�[/]T�,E6yJҋ���(V,���(��a_�ς%������Iڼ��N�Ը��ϯ��ş
1&��H<��#�&i�	�K�&%�I���d�k�q�A����}�����٪��;��>1��� &�/;��L��t�M +e�@����V�1E�*�x�>TZ`��-�h��E޻k�9�3�p���������#�T 콆��]?xc_�4X��2�{'ml�3!��.u9�����M����#
��ٚ�}���^-Q2��K��;�����y�D��>�W�k���s�����$�	5�ȟ�d6w�̇�6ʔ9x�nhv#�gm�C��*�>p*�̐RN�
ya]uԺa<	޾�&�	7/�!Q���>p\u���b�(F���2�����o0�yф����恘�U9A�|�~uB�������Ӵ�*+�f�j�K���
�$�f��ZR<�M<�J��Ǔ �U<;���(���q|��*���K��^aZ��Ǳ�Ǉ'ȹ�c��g�`n�7bP7ż���.���n��.e��������Ek۬�V�xi*��?����;Vq���#J=�m�������9P1�"^�ٕ��ckX~�ֵ�-�h����u5w�_�u��x��&��-�>�	�b�s��s�^@k9mIf��2i����1������_<�|�
�̻�.���/"N=z��Ti�s�?����jr��8�z��eW����̑���G	�}$�ʹĻ�!/�<!?���cZ��W�����s���շ��zC���C�����7LX'4��#���O~���Z1�>Exc��C�� Mk� ����z�������B���8W3���s���Y���q�1 2@��TC�2��#����փ��` e f �w�W� @�w��f��q?G�^ ����'�L�;�%�ߋ���v��ꋻ���ծ�K���c�5]/�J� �M�^�AxZ��A���$Z��X݅��X\W�+pδ���sCiE