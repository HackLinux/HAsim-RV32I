�
�t��#��4ƒ��,����Y(f�d�	7�MS�e�b�T+!�3+-i)�Y���B{;<v�Ñ�w�e"9K��($$i������Dl� ��7�q}.	 ��x<"��i���ƕ�L��0�R�ҭH�Sp��L�y\7Rv�7(��߭:� ?�$�;�o��+����%��ZS)�p�d
�z�������,;g�.�:�o��N&Ĭ��m��c݅�Z�\� �J���
���)h
������Lt$����u�!"@�U�+��ڇI�w�&�u���+�3���j���lf��B;$GL
sY�����\;��}��p}0���&�!�~���w�U��������gͱ��v�v�I�R�6G�5�������*B��Y��d��Κ����E�IІF6N�1>�z��x&���j���p�'�f���A:�p0h�P7:�G)|� ,��c�v��<�J��b&!+8l�����NsrH��?Fv��
A��F�����Y+8�nSj�(ӂ��d���������v�1��굻�����nrE�1���	j2�-�oD�����T����Dם�{�fR�I꠪���'���ԃ�3�$@����:�̏ba���fWg�R&�j�a�V�lô~Y\�gx(t��^`[t�g��g��_d��Ј�ۨK���G�8ǥ��u��^��M��R�[�:$�x~_���r���4�䀧�,���8� ��ɝ5s��-���Q����\z��EC���8�uS>	�,,��Ò�R� l=���i8���n��x�<��4�-�˰R��K����f���<��֢d��u�H��@���	�_N~�sߒ�,|\ $ZV��k��v�-dg�T�a��$M��$�	�~�Ç���J�? ��|Hѡ%[��2��+o0�J�
w��8w��-��-���Pb�
�G��=�$����1a�Ӡk�P���C~u���o�G��mt������Cd��"�K�T�}�=��"C�a�$畠q�fB��`�d-X��Z>�)e�ݹ�7c���C5�U/|����*�$���AKӝS��D���τ7�}(�Ui(��
&p��}�D2�Er[�8A��uz�(p��xZH�-��gQ2~Oߎh�ݖ�;6@`��(hA�;fJ�R}=����T�ǿ�D�^��1�}�}�Я��實h�_�}�ZA}�`�yY&>+�}l<6����|������ھ�}�7�Dy���8gy@�e4��!o�N�I"�"Cؘ��EjY���dE8���� �,��xlE�u�򶦛`�a�eU��X���0޲�1�ank�o���r�.}+<m�:�-~�J�X�Rv!���Da�I�4Q�O��W��77��N� ���T�3g�=RF4a�Kq�X:�"�aB�a�IB������1��R�Ɖ���@��3�1�J��t~�Q��,��O+kD�/��uN]#$�����_�=[�z�q�������n�5�A�4
������68����a�J�{1�v7�6���7JcY�B����<�``q'�:BҝS(��L8�I$6!��Z��X<��~�`�{C�d��o��[�Uj]'����ޖ�~�g��X3����q]c��/pw�8�������������t/>d�4E�u��H~�IX��6��1�YN��Z����4�����޽Ql��˹�gom��(Y
�?����s*J�"�x)v1�_�OA��rj�8����7yfO��s�ŸO��#f�:z\������sS���8X��ij��Tb���:�A`���J����#`G�ݻ���[dˇ��2�͚���g��3&K^r�/���y����P�������enޙ� Y$Eg8�� ��%�e������ҪU���ciE�"�.�@��Id���?���f��!��_�rm<�Y,��<��'g��\b�B�ͤ���X]���>%����0���B�8�?���cD?�C�V�)�W��P��I�����<0~��a�Fotz�K��@��Ӏ�^�E��sٓ �<�gʤb���q�y)�z��1��p!�-��a�
$������~�|��q�d��H;�D��h��&�[�<99.k��+�ɑ֜ڂ��|�������pFk�z�O�C4�[� �Ŝ/ى��c�C�q�c�/���e��;6	F ��P�x�lX�㥏$��#WX�#[	�|�zТ���a1�m���楎õ�)�����=��p�8&Gϟm/���Ͻ�\���L��\w�y����ʔ���R�� |�i,��a`�~i�8���N]���*\%�� `���l j9���Y}k����A�iN��>�M��/*6E�&A�&�ߥ+R۱�$�1�5���b��qGyČ�+7m�W*a`YG}�`�����/�C!�J3��~��YiUL�>Y�e�"g$�����`�q����j�U-#��ȅc�g	�y:s�0�k���Z�=�6�c!�%�@%]q�ض��1���4�&Y ]��r�7��2��O�IES����3+5\�:	Nx;,�x5h��t���)�C�e�+gAחE
�r)x�л����-��!�1���|��>�z��{�/�`�_/��#�|�I���$6{ښa�E��Hd1��e�f��a��`��	�H��/��3��B�4\���q~	�F���g�2zΰ���gɏ<��t`�����})��۔8���\��UY5A �d�{�.���Y�7�U�z�V�����-�V�0�ݰn��|r���}Q��h�ӡFT����Ӵ�G�(5]?mz[Z�e�����S��fܗ�w)�J�d���%��#�E7,�B�O	VD@���ƽr'y
P3� �_����
�;$���Q���~)�~4�*y�r��-ZI�FLP�0 �#Rv�o���GAQ�8����'#�̭������_T�y����<��R*қ��Ls��ӓ�ڨ�݋l�m ��ԏ6�6����/�ɯ�*�Y���/+ 4���@F����Y�o!]�$^5ov` ������￥�lK��V�ێ!�������ʽO����G2B�q�=׼��L������������JF4^u�Ȩ��=� �T�U^��?�z�M���+�Kp���Kt^�ӎ���߿Z�/C�Q���۠�O�ٍ��G��(hT`�lU��ـ�a��k#�S����U�v�CƁ��ާ��P��_�҄;l&h�8n*����N�qX����dc~Mvz��n�ҕ3$|d��ιp��}N����G�M��?���s�Y��# �ޜ}�����hԜ�}����mʗTT$��k�)o����xj�į~�=��M��Q��Vl s���ƿ�y;�]q��HK�2qطN�Y��mo�8�ⅵ��7��.r��T��[2�*�h�['��깿I�ĥ��괮��l��m#������A��v0?�˦�����J`�i�3��u��S*����o]���d-#�el��ѷQ�4�	�Je��%0�h��j�}�j�����_j�M���������Yoh3��5��K�c
�cng
�^�f�S�+�Co���7�'sq��0�����VX�aW���EG����FZ%��m�&g,$d�0���li0:hR��s�M|��CbY���B�I���%4�/Ƅ�kp�e�T�#�lq�d�U�"a�(�d>���j'�H�~r��w嬨�e�+�B�lmWf~vB���>��!ˀ/�DF�b�%��6�(�����a�c�Q��'b�z��VYl�G�B����#t���� ��o�Y�)�w^��M�Ό��T �0�&���w�&a�m��-w�'�g���ts���w
�N����P�:����f���j�9�D��i���5�P��s"1[�=}AL��?��J��������]������G�v����w���v����m�y�ų(��q/��'����������r�j��j-����5�b/r�E�0 �G�u�rƺ�����"-q���۰�#b4��� �1C�������a0���% M���pɯ@�`����j#�`��SM�/S<R���z���5�+D-�+O�K�4��Z���x����s�G��@FN��m�0 �:H�hS���=�}S���1R�x���|X[4s*�F����XU,?�N8\���̌�5��6��c�t^m�
p�ÿF�w�2���񮞚��p>��{i׌��kG�fa�5%�ܓ�)P��qP���Ib�U�5�y/r�BR:<��:��O�~�C��c�|�.��]�|�h�K�8�I������v�\�cj�Y��}]4q�!�S��0�c������rA�Hu���0T��WgĴ��`�n���Y�x������a�F�{�+x�vp���\��ww��B�������C�~�u�#�ɭ�M�C��ŀ�RxZI��,Q3�m)��3�+5�Q�j5��'FXr�����?�����L�G@Ї�g�Ţ���+�v*�<�G \��g<�I��� L��
����O�b�$�Y�W_nKs,�������a�����z�s�joSK8G�N5q��has�)���,o��傒(M��<#�pʨ�h]��ɢ�p �*��b�u���4x+�uz�Z-��Q�M���+��ȕP�E�0_��ݛ����QqYHm�U�Yʹ�)���&v�U��S>q8��RZ�Y�Rľ�k�`Һ�>&b���c�2���B>��q�ra��[��B�#Pҡ,v�F�M��+w�v�\�ss��帗!2��
 %������5`e�i'�GL�M0��9̩!�ެ�$S!5�l�;e�����9�+�*�T^`{�,�T�͋z�I�M�ÂH����i�\���u�2#��D�O�ė���q��C�O��3%���um��p�[j�+,�W/��="`�pyMRVo|�^4j�6���7B�8�.L����^����5F���"���S��L���M�{ ŧ"ؠ��r��	c/�r�ю�NA0L��1P1���[��U�����`�����ND�,�����Hr꒴�!�����0��f���`aG��^F������)q����������InEy�YK�p`D4�K��4W��	������x�OE7#�ᯎ��=H�W�3	:Q~�O#��K��F1[�Ј�o9QI�H����<	�� �iND�?���m ���c#H��K���~��p4H�0(WM�4X����1����=����Ȟ#�������dI�7�����'�$��R7{���Wd@�~.��~߅���s��xnw8�a�1�C�@0P���|�1�I���Es(��~�O�1�a@	Jv�6~�>H<}�]�TC�R�p���9{�y�=nH�X"jB�E�h�#�9P�L��!T����vג ��LL�۶�Y�&�����f��M6=��۶�ER�U/V�T�"w�P�>���?�h��/#�s��<��G|t�ݤ-cZۇŶ&߆I5��D�3�)>�n�	炶0[%��x�b���N��`"��7�8L�$$�^��BV�c\�1Ou4h�!G������t��"��W�p�?��u��:n������Տ�� �[�+
�B�Q��H~���I#c޾Nx�WE7'�ėB6N��Ԣ#�A��ֈ�S��	�Ყ����爻4<g"�1���`T�^Ca}�c�,o��|g��)�[�c$;���7-�]��ߎ�3ADaz�0M+J*և�q��!x&͢1��M�	���	���Ui�+�:W������3:������ℍ2Җ���I��#�=���Ő��#�Q�ϯ�����O�꓿u�h���m�b��Y�;@��@��<T`�/p������b�INA�k�
���ۨӌ� \��N� ��(Z+�𾣨E�tiWn	
dj����n=��9�ǉ��G:�(Ӣ?f�U���gCy�1��(�A�����k��Dc�O39P2�?�բ�@'��i���1K:��҉��vfG���!�:�ֈ��+o�IE/C�T�e�y�V���7Pz�#����T�?�vPc�#M4m�6�;V�� %�b�T9���V��A�JDh��N��`��)E��2�c�E~�6��1��p��^���һcה��F�m�Or�'�T:n�Ux���U�3f�_�x�M��RlcTl��$���|S�j�U�XI�İ��Ov�����0�(��YΠb_��A�
Iw]ڴ��#�N{�m�^�FEY���1�N֬A�.��;yc�6��x���I�_�pK�{�]��3��r{�!�:.��̝$�~�M��������&S�U�r$"<ӛ��ػ�{,��������$�i�av�~7P�Sn�g�T8Aq��*�Cz�rS�*�tJƫh�dȆp���|�m���Fg'��1LC+�{�m�$�M��/}ɜ�dA�duw'�vB~V}P^@�bU�o�Ʀy�Pg@�M
�@Dw'I+�GPxHԗI�v?���Q�ո�����\1�V��U*�6����:��p)�7�$���Le�$De�+Ko��Mz��Q}K"�D���C�&Mar�hǾC�D��U�٪�g
{B�x��J?U�Q���*r|z�Y��OA�jJ=\@ܢV�{��.�:x"i�I.#�NR׏��/o
4�V����o��}���3$��@��z�����}r�T{��N+�AZV�����P�"��=��5�JKL!�$٨g������'����ӎ\*�A��A"G�xc������%�[���i��	�:=`�&�8؊CT������`p�Y^��������#����ml�z�8��2#�K�v��v?I�O�j)�m�3$�U��	��?U������]�T{#%"�:U���0-�,�ғ���6��|�^�����6��I��b����týu��H:��;"���8�%�)c��So�DΜ�:��Q�_������%ҸR��mE����N�G�[��&��߼c.�<���AW�f��]�����&J(����[�X`��Ϭ��I��EYVZ�
j�k<�1��Tt��]U���J�r|�-ŷ���O�ig?�a۾M݉l 6�� wa���2**�4/YOإkĨK3�hVoK��d��H��X�c��I��QS�k���b�T��,Ja�zE�I�Kf���K�ֿx�Gd�������D>DI��S6s�Q��.�ry�	`���ZD����8EV�x����c.?��X}��ú���9S��o��x2�FY�z z�r��� ��I��=u��e&v�-������t��Zݡ ���꾗�|ϥD�~`^�����{`��J}��@\_'z����y����c!��^J*�3�%��7-����^��Bquѻ��آ��!��q�[� ��0(�ш�D*������80:���A�Q(f�E�������Q�����2ͤIË	�