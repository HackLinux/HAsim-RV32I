������ﶟ�����������������������������ȝ����������������»�������������a���l�������|ߎ��Ŏ�ŋ������u���!!�!����!���������������������ǧ����������������������������ŖŖ��t��!��y�y�y���!��궐쑐���������������������������!�!�!y�y��!놆���꟟������������������������������������������ȝ�ڤ��������ڣ����������������ˋ��������������ߋ�ߋߋߞ�������u�q���!!!!���➻�����������ǧ�����������������������������ŋŋ���������st������[�[�y��!��u�������������������������uu����!�������!!놆���u��������������������������������ȝȝ������ڣڤڤڤ��ڤ���������������M�M��������ۂ��|�|�|���߂߂��u������!�����ꄒ�������ʧʇ�������������������������������ŋ��t�t�ts���������y�y�y��!Ά궶������������������������uu��q����������!�!�q���ꐐ��������������Ȑ��������������������������ȝ�����������ڤ��������������ڎڣڤ��MMMM?����������ۂ���߂��߂߂����������!��|����������������������������������s��s��������s�t���s�s��!���}�}���!�궶u��������������������uuu�q�q!!��y�����!�q��궶�������������������������������������������Ȕ��������������ڣڤ��������������������MeMe�������������悂�ۂ�߂߂���q����q�q!��⋻�����������������������������s���������������s�s�t�s�st�u���y�}�y�熆�궶u��쑐����������u����ꆆ��!����������!�궶��uꐐ�ȑ����ȝȐ�������������������������������ȔȔ����������������ڣڤ���������|��������lLMeM�l��������������ۂ����������������q�!lqX�������������������������������������������������s�s�s��u�������y��!�q궶�uu�u�u������u�u��q�q�!!�����������!�q���u�u������������ȑ�Ȑ�ȝ������������������������ȼ����������������������ڤ����������������~�aeMe���������������₂�ۂ����u�������q��q!l�v�����������������������s��������������������������t��t�u����������!�!��q궶��u�u����u��qq�q���������������!����궶����������������Ȑ���ȝ�������������������������Ⱦ��������������ڿڿ���������ڤ���σ��|�������aMeM����l�l�������������ۂ삂���q����q��q�33փ�s������������������������������������������tmm��������y���!!�놆�q궆�qq�q�q�q!!��y��������������!��q��u�uu�����������������쐟�����Ȕ����ȗ��������������Ⱦ������������ڣ������������������ڎ�|ߤ���¤���MMMM?�����l���������悂����������q�������l�|����������������������������������|m|��!}�����������!!!!!������!!!!����������������������ㆆq�u����������������������ȝ�����ȝ���������������������������������������������������������ߤ|������MMMMM���L��l�����������߂���������q�����!��u|���������s�������������������s��u�����������y������!������������}�}�}��C�C�����������q��uu���������������������������������ȝ�����ȟ�������������������������ڿڿڿ������������������ߤ����P�������L���l����������߂�������������uu���!q�������������������������m�|m�����������������������������}�}�}�����������������q��uuu�����������������������������������������ȟ������������������������ڿڿڿڿ���������������������������������������������ߝ�������������������lqu�|��������������������msmmmq�������������������������������������C������������qq�uuu����������t�t��������������������������������������Ⱦ����������������ڿڿ����������������������������P�P������������������������ߞ�ߝ����������!�l�|���������������mmmu�������������������������������C�������C�����������q��uuu�������t��t�������������������������������Ȑ��������󗼼����������������������������������������������l�W�W��������L���l����������ߞ��ߞ���������u�����lu�����������������mm�q�C�6�6���6�6�6�6�6����������������C��C��������l�qq�uu�u���������������������������������������ȝ���ȟ���������������������������������������������������ˤ��W���W������������������������ߞ�����������u�������||�|�������������ms�����6�C���6�6�6�6��66�6��C6��C��C��C6�6C���������q���uu�����������������������������������������������ȟ���������������������������������������������������������WW�W�������������������������ߞߞ���������������⃃����������������m�u�\6�6�6�6�6�6�666666�66C�C6�6C�C6���C�C����������uuuu�������������������������������������������ȝ�����������������������������������������������������������W�����W����������Q������������ߞ���������߂����������|���������������mmuu��C6�6�6�6��6��6�6��66��6�C�������������C�3qqquuuuu�|�|���������������������������������������������������������������������������������������������������������������W��������������������������������߂��������C��|����������������mmm�uq��6�6�6�66�666�6�6�6����������������l�q��uu���||��������������������ߋ������������������ȝȺ������������Ⱦ������������������������������������������������Q������W�W��������������������ߞ����������ߞ߂��u������l�~�����������������m|�A�CC�C�6�6�6����6�6�6����C��C���?�333�qquuuu�||||������������|��������������������������������������������������������ȼ��������������������������������Q��P�P����������������������������������ƺ���ߞ�����������₃�������������������������|muq�C�C�C�6�6�6�666C�6�C�C��?C����������C3�l�q��uuv�|||||���������|���|�����ߋ�����������ƝƝ������Ⱥ�ȗ�����������Ⱥ������������ȝ�������������������������������{��P�P�P�P�P��������������������������������ƞ�����������l��ゃ�����������������������|vu��}}}}�C�C�C�CCCCCC�C�C?C�����C�C�C��?�����q��uvu�||||��������������|�|�ߋߋߞ��������������������Ⱥ�����������������Ⱥ���������ȝ���������������������������������P�P�P�P�P�P�P�P�������������������������Ŗ���ƞ�������������⃃����������������������������X�\�}}C}}}C�C�CCCCCCCC�C�C�C�C�CC�CCCC���l����u�X���||�|�������������|�ߋߋߞߞ���ƞ��������ƺ���Ⱥ�������������������������������Ȕ����������������������ʻ������W�P�P�P�P�P�P�P���P����������������Ŗ�������ƞŞƞ�߂���l��aւ���������������������������v�A3����C}C}CCCCCCCCCCCCCC�CCCC��C����L�l�������u��||��|�|�|�����|���ߋߋ|������������Ɲ�������������Ⱥ���������������������������Ȕ�����������������������������l�P�P�P�P�P�P�P�P�P����������������������������Şƞ����߂�����l��l�~�������~�����������������v�q3���C�CC�C6C6�CCCC�CCCCCCCC���C�33�ll�����u��~�����������|�|�||||�|ߞ����ߞߞ����ߞ����ߝ��������ȝ����������������������������ȝ�����������������������ʻ���QQa�Q���WW�P�P�P�P�P�P�P�����������������������Ş���ߋߞ�߂����������l���������~ۉ������������ۃ��L��C�C����3�3���CCCCCC���������all���������X���������|�|�|�||�|������ߞߞߞߞ��ߞߞ�����������ȝ���Ⱥ�����������������������ȼ��������������������������»llQQQQQ�����P�P�P�P�P�P����������������������������ŋŋ����߂߂������l���l~��������~�����������������L�������qqAqq+l\LL�C�?�L�3�3�3�l���������~�ۃ���|�|||�||��|�||�������ߞߞߞߞߞߞ�Ɲ��Ɲƺ����������������������������������������������������˻ڻ���QaQQQQ�llQ�Q�W�P�P�PP��P�P�P����������������������������ŋ���߂���u�������}�l���A��~�ω������������~�L��d3l$�~v���v�~��(la��3�\lllll+���A�����~�ۂ������|�|�|߃�߂�������ߞߞߞߞ��ߞߞ�Ɲƺƺƺ��ƺ���캝������������������ȼ�����������˿������������Ƀۃ��Q�QNaal�����l�ll�Q�QPPPPPPPWP�P�P�P����l������������������ߋ�߂�������q�l����������⃃����������������d�*;v�����������A���3l�������q���������v�ۂ���|�߂߂߂��߂�����ߞ��ߞ��ߞ���ƺ����Ɲƺ�ߺ��캝������������������͖������������������˻�ˎ����NQQN�Q�l�l���������llQQQQ��WWPPPWP�P�P�P��������ߋ�����������ŋ�|�߂���������l���}�����l~v�����������~<lda�v�����������~���l����+l�+�������������悂��삂߂߂������������ߝ�ߞ�ƺ������ƺ����ߝ�읝����캝���ȝ�����������͜͜�����v�~~���~���~��{�~FFNFQQNl������������������llllQF�PWPP����P�����������ߤ������ߋ�߂�ۂ��������!l���e����l�~~ۃ��ωω~��L?C�3�~����ۃۃۃۃ~����a�(l�L��ll������������������������������ߝ����ߝ��������������������ߝ��ߝ�ߺ����������������Ⱦ��������͛͜�.ll'(��?��'a%WWW�F�Qaa�l��������~��������������lWWWPWP�PW���������ۂ�ߤ����Ŏ�ŋ�ߋߞ�����������l��ee�e������ۉۃ~l����L��;~~~�~�~~~~~~~~�DlL����L��a�lllll��������������������������᝞�ƺ���������������ߞ������������ƺƺ���������ȗ�����������͛C�^)kk))���dddd&&�W�F�ccl��D���~�~�~~�~~~~�~~~�~��laPWPWPWPWPWWQl�����ߤ����������������������������������������e��l������_�������~�~~~~{~�~~~����[����������������lll���������������읝�ߞ����������������������ƞߞ�ƞ�������Ƣ��������������ȗ��������������O^k^)kkk)k))��ddd&&�''����D�;�{�~~~~�����������~��aPPWWPWPWWWWQ�����ߣ����������������������������������e��[e��_�_����Q��{~{~{~~{�{�{~����L�e������������������������������������������������������������������������ƢƢƢƢ�������������������������kkkkkk)k)k)k�)�)d)d??FFa'����B�{�~{{{~~�����������{~��FWPWW�WWWWQQl�������»����������������������������������e�ee[e[e[e[ee�l���{���{{�{�{������yee�y�����������������������������������������������������������������������ƢƢƢ�����������������������������kkkkkkk�k�k)k)kd)d�d&?FF����;{{{{{~{ύ�����ω���~~��7�iPiPWWWPWPa����ۋ���������������������������������������������e�����������������������e}e}�}��������������������������������������ߞ������������������������ƖƢƢƢ����������������������������������kkkkj_j_jjjddjd�dkj)dddLL%��D�;{~~~{~{ۍ��������ύ�{{�G��PiPiP�PWWQl������������������������������������������������������������������������e[e}e}e}�e����������������������������������������ߞ�ƞƞ�ƢƢƢƢƖƖƖƖ���������������������������������������jjjjjjjjjjjjjjjdjjjjjdd&d&?FQ'��{~~~~~~~�~��������ύ~~{�cNiZiPPPWWiQQ���ۋ�����������������������������������������������������������������ee_e�e[e�eee}e��e����������l��l��������������������ߞ������Ƣ���������ƢŖ������������������������������������������jjjjjjjjjjjj�j�j�j�j�j�j�jZZ&WQc�84B{{{{~��~�~��ύ���{{{��c&�PWPWPWWWW���~ۤ���»����������������������������������������������������������ee_e___e[e�__e[e}ee�eee�M������������lll�����������읝Ɲ�ƢƢ����������������������������������������������������jjjjj�j�j�j�j�j�j�j�j��������WQcG:�7B{{����ύύ�~~~~{{�{���WZZZWZWWWWWQl�����|�ڻ������������������������������������������������������l�ee�_e_e_e_�_�_�___�_�QaQaQaQa�llaa���a��a��ll������쑝�����Ƣ�������͕͢͢͢�������������������������������Ȕ��������jj�j�j�j�j�j�j�j�j����idiii�YY�GV��7�{�{�������~~{���D��D��QZZ&Z&&WWWWQ������ۃ��������������������¤����������������������������������Q�Meeeee�e_�_����QQal���{{{~~~{~Ϡ����~�~���l����l���u��쑝����������������͖��������������������������������������������Zijijijijij�j�j�j�j�ZiZii�WpN��VG��4B{{{�����~{{{{����0��ldid�ZZZ&&&Fl(������~ۃ���|ۤ�����ڎڤ������{���������{{�{{{�{��������{���Q�eeeeeee_eM�Q��~����������Ϡ�����������������~~�l�a����u삂���t�t���������������������������������������������������������ijijijijijijijijijiZZPiP��QQ�p���G����BB{{{{{{BB004%%��D�%adddddddddddd&LLlll+���$�~~~~~��ω������~�~~��Ql��������4��{�{{{{{{{����a&�j_�__��Q��7�~����������Ϡ�������������������������A���q�u���tttt����������������������������������������������������������ZijiZijiZidiZijiZiZiPWW��NQ�p�����8�����00�440004/f%8ff�'adddd�d)d)d)dd??La\**DD.D;D;2{�22{;2~~{~���aFQa�l%�����04�4{�{�B00��Q?___j_d?'�~~���ω�������������������������ɣ�˻�ɩ�����X�qq�u�|��ttt�t��������������������������Ǆ���������������������������iZiZZiiZiZiiZ��P�W�W��QQQQaQcac��������88���%%�f%%'aj)d�ddd�d)d)�)�"6�3l\�+((.(.( (��� D %�%'aFLFQc�8��00B�2BB�0D�%W�dMFG/02~ω���������������������������������������������|v~u�uu��|���t�tt���ŖŖ���������������������������������������������W�W�����i������YNaNacQaaQQQQNQaQQaa�������%l%\��*��aa6)d)d)))))))�)""�5��  � q +((++**\aaaaaQFFF??FQ%%8D�0�B,2,�D%a''B~ω������������������������������������ɩ����������������|��uX��|��������t�s������������������������������������������»���������Ncccc''a�llaaca�FFQaaaaaa''�aaaaaa�aaa\3\33���))))))))))""����qq�AqAqAqq+�\\\33L???C???M&a'�0,�;�;0��~����������������������������������������������������������˻�����u���|�����������s���������������������������������������������NN���NNcc�c��%��*�*�+�((\�l*l�lll�lllllaa�33a33L33L���C"�)))))�)�)"����qAuuuXXuXX�$$A�+\\3�CC��)dkdk�k�k�kjk?Fc�%8��D-��������������Ϡ��ϠϠϠϠ����ϣ�������ɽ����������������ɩ�����ˣ||����������������������������������������������������������cNN�NNNN%%��%�����.D$������uX�u�A�Aq��llllaaaaLLL�LC��)k)))�)))))6�\�qqqAu�XXXvXXXX�$$..+*\3�C�k�k�k�k�kjk�kjk��?Fac�%�D2���������������Ϡ��������ϠϠ��Ͻ�����������������������������������������������||������������������������ˣˣˣˣˣˣ�ڻ�ˎˣ������a�a��������q�A���v����|�����|������v₂�ۃ��D ��F��)kkk)k��C���))C3\*.$A<<<XXXXXXX~<<<<�$;D(%aF��d?�c8???��kdk��??F'D�2~���Ϡ������������ϠϠϠϽϠ�������������������������������������������ɩ���~�ۃ���|��������������������������������������������l�llll���������잞��Œ����ʒ�»�������ɻ�ˣ����ύ~�;��L�3LLLL�L��}}L\��D;;#<~~~<<~<~~~~~~<~~~$;�(�aa'%;B������������BB�{����Ѝ�Ͻ����������������Ϡ��Ͻ�������ɽ�������������������������������������������₂���ߞߞ�������ŋ������������ŋ�tŋ����t������t�����l������������͛�ǛǛ������ˣ�������������v~��\�llll�a\�\���\�.�$$#{<2<~~#~~~~~~~~~~<�9;D�(�;~����v�����������������������������������������Р�ϽϽ���������������������������������������������������ȝ����������ƢƢƖƖŖŖŖ����������������������������������잞�����������s�����|����vvvvvv~v~v~~~~~~(�\+�+�+��ll\a\l��;$~�~�~{~�~�~~~~~�~�{;;��*�09��ύ���������������������������������������������ύЍ�Ϡ�������������������������������������������������������������������������������������������������������������qq�uu��||�������|||m|mvvvv~~~v~~~~~~9~2#;;D\a�l(�(+�l*a\al\��;��2~2~{~{~~~~~{~{~{{;2�D�{�����ύύύύ������������������������������������������ύϠ������������������������������������������������������������������������������������Ï���������������������!�qqA<XXv~v~���������|�����������~v~~~~~~$-�ll���������laaal���2;{�{�~�~�~�~�~�~~~�{�;������Ͻ��ϽϽ�����������������������ύ��ύ�ύ�����ύ�����Ϡ�������������������������������������������������������������������������������������������������������������  $u$X~~vXvvvv���������������������~~����.��.�D.D0DD��l������~{~~~~~~~�~~~~~~~�����~������������Ͽппп�������������������Ϡ�Ϥ��ωω����������������������������������������������������������������������������������������������������������������!�β�����uXXXXX~~~~~�~vv����������˻�����¤���~��~~~~~�~�~��$����A�~ۃ���||�|������|��������Ϡ��������Ͽ����������������������ϠϤ�����������������������Ť��������ǖǒ���Ǜ�������������������������������������������������������������������������������!!!���u���������v�XvXv~v~v~v~vvv�������ˎ��||�ߋ�ێ��������������₋���������������ŋ�����⤤��������������ڿ����ϿϿп���������������������ʧʧʧ����������͖͖�Œ���������ǒ��������������������������������������������������������������������������������������u���������������vvvvvv<X~~~~~~~v~~~~~~~~�����������������||||��s�������������������ߋ������������������������������������������������������ʧ�ʧʧ��������ǛǛ�ǒ�������������������ʧ��ʧʧ�����������������������������������������������������������������u����������w���s�s��������vvvvvv~~<$.$<~~~�vω�����������������������ʛ�ʛǛ������Ȑ�Ɩ�ʧ�����������������������������������������������������������������ǒ�������������������������������������������������������������������������������������������u���������������������������w�wmmmm��uu�mm�mm�������������ω�������ʧ����������������������î����������������������������������������������������������̧�������ǧʧ��Ǜ�ǒ����������������������������������������������������������������������������������XXXv�v���m�m�w�w�s���m�����mmmvu�u�uX�m��������������»»���tt���������������������������������������������������������������������������������������î��������ǛǛ���������s������������������������Ŗ�Ɲ�����Ɩ��͜����������������������������������~~~~�~�~�~v~v~�ω��ۃ~~~~~~�$.��.;9~~~~~�~v������������|�|�����u�|���t�������������������������������������������������������������������������������ç���ʧ��������Ϥ��������������ω���s�������������������������������������������������������������������mmmm�v�v�������~�~~~~~��������<~~~~~~<~~~~~~~~�~v~vvv~XXXXX<Xuu$uu�u��mwsssssstmwwu�mr�������������������������������������������������˿��˻�����ʻʇ����������������̇������̏̏����������������