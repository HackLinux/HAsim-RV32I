�a3b4SbFvbT~bJ�b4�bL�bU�bGgcN�cL6eKQeG�eF�eHf;/f"0fb�fU�fB�fJ gB	g5eg2�kB�k;8l>�lD;mLgqG1r3urLsU�sB�sGt=(u6;uLYuI�uQ�v4w9w4�w+�zJ{O,{?I{J�{G�~;�ǸQ܀K�H��P��GňQ��C��H��=��.��O��U�@b�7p�DߍF�Q{�Pُ=ۏJ�F��@j�+�E(�C6�PC�I$ �[�_�vǏ,��%`ObN$4Y(WO�
��:N;N�Y,1\!�a*/f%s/�w$��*K�$(uV��b$`O @T1PT3JUb'�� N#	�*N�N3b
�p*�*p�)�&�e ��Wɋ�&$a�$(;N	`O5�SBb6�v�>�DǏ1m�6�+Yu{�%wP"T)�b&�v%p��$0R!�*<�
�N(`Ob��� N2;NA�N;NO<P?�Q80R*�R&`S<�S3�S?�V6�Y?\A _,�_?Sb8~b7c?�cC�c3>e2eg9{k-rB,r?1r6t2(wCaw<�w4�y0�~?ɉ9��*�#�1p�4l�<��4 �Bw�GU�B'T'�$�N�^!b�g'�$#�`O"�_
b$�l`Ob;m[r!�v�"�& N$wP<�S0�S+5T8�T1�`<~b3�b8�c2be&eg.(u4�~*��.�ߍ&�5�vP�:׋1��5�[V{ o`OY��;N6�N8�N&VS'�S eg!k?�s(�v�~.D�(���*�.b�7�N
 _ Kb#pe%�{'Mblx ��v��(u��^Ǐ�[ ��v��kN�:Y�w_Nb$5ub�v$�_+a-b$Kb0�.�be_�[Y�_�$
N O!�O#HQ#nc	g�(�[ �[ � 3$>PGRD@T@JU+�UG.^8r^?S_>�aGSb8�b9�c;9e6w�{?�~>ɋE�.�1Ǐ*��?��:�1�RN):N=O$OEUOE<PG�S?�S4(W&\@�`:�`L?a4�a3�b>be6fE/f"SfR	g0eg;�kG1rEtGwAw/�w�~<��M����<��7�@�4�Jj�I�G$�:(�7�[?e fck*N*�O5�Q0b1%c%feg;�l2kp8�s�v�w2�~2>�9"�8w�1Ǐ7��?�2�N�m܀$O.�v(�vZ?�E�b��/f���N3�NC�N$`O�O9vPC�T(yY1�[1S_Ib/fF�gF�C�/�?=�Wُ5��<��F�N�OC>PF�RKJTF`1mF1r8�wB��/$�N!0R/JU1�c/�v�#Ǐm� ��2�/\O�$�S+PW%�` ab#w(A��`b�$�'$ $$`O-0R#JU0b+�lD�v��+��.Ǐ�)�%�,b�gb$�8+R5b8}v8ɋ $$ �N`O"�O=vPER=yY:\=b���.$b�$jx$$�T$$!k
�S�l$&;N2Lk�v
�-Ǐ-�� ?$`O4b3/fEwE�8ُ8$b�"k $Y�v�!Ǐ��!��5�${ �] _ Y�[eg�(:N	1r�!� C$0 NNN	NCNCNA:ND;NJNN*pNN\OL`O0ZP:wP=�PTsQ@6R-MRHVSL�SZ�SN�SUTA,TK@TQ|TK�TI�TU�T7�TK1U;JUCY?YG'Y?)Y?f[B�[S.^Lr^Kt^?^B�_D�_F`Q`I�`L�`3�`Ua<b(SbCnbP�bQ�bMcPccR�cO�cPdG�dU�dS�dQ�dJ>eCceQreF�fBmgH�hB:kPlQ�mN�mQ1rBurO�s:(u6{vJ�vUw44xP�yL�zJI{:�{M�~N�~>�~A3�L̀>9�Q��@ŋU�0�<ߍC��<ُ/܏L��M�U �N��6D�AL�Qj�EΘI��C�J�L$
�!$;N#(W�^�,�cUSl�
Xdt	�W;m N�S2T$�p&�#�)N
��b$JS �T%�U-f[#�["Zf%n'7r#ɉ-�)YuQ�'�R�SK`g w
N'Y�N�Q�Y$ N,N2�P-JU4�Y:�[71\+�_"b7Oc?Il:w'��:���:��-�)�$7�??a"�g
dk0Rb�`O�7u(WP[ `N�v�&Ǐ)�$7�pa�cˆ�vyb`{k�v�#�$"N?"NE_N@pNJ�NHPMZP:?QF{Q:�RHTD�TS(W5'Y?sY;�Y9i[-\,\L1\Dt^J>eI�eA	g �nAvpD�pJ�rE�sK�v�~I�J�?��AňG��>�Np�EُE�NG�I��5��9̑7�A��Jb�; �K�>�K(�6K�<f�[ eg�v&�#�$$N$�N/`O!yY;b1r@�rI�2��I�
ُ5{k	o�|	;N6�N6O%eQ=�Q+�S6:Y1\B_2�_Bbb6�b:�c.Xd7/fKf> g.GoC�p>�p={v9�y;{>܀:��$b�2ۏ-�8$�e�r!�,�
NBN)�NKO HQ:`S?�S=�SI�SB�S)�TI(W9YK\1�^?S_@�_:`RSb8~bF�b?�b.�c2�c?�eH/f gA	g){kE�lG;m/1rB(u9-uM�~B����;��=��0�D%�Mb�/ߍC��)��H�F�8(�;B�<�s�v$�n \O�S�ZW$�~$gU
OW1�Y4b�v%p�"�-7�%`O!.^(�_b�~=�9Ǐ<$JU/;m.�n8�v	�'Ǐ*�$\{�N���yЏ�[{k/ɋ&��$���$�S�Y!�g4o7�v�4f�-n�<�+b"N�v�$$xY��$%;N2uQ*�[$�[(9\=;`3b,?e/g0Cg$w	���/��8�T bb�P6�{-N o`7�`$t(�u�u(�x'o�,̑{��_�!N�$�z$�S&eg�p!�)}^!�l!��`U[��0�$�~$JU.<w.�b)/f�~1rb�\Od�` 1Y�N?a�us�	�v	 N5pN7�Q0R$�S$�S?�S8T(,T6�T41U=�U:(W6b(�b96e=eg.�v/w+�w7��Ջ?�Dߍ2Ǐ,��D�8`O%`1�`5b�v)��/7�5tQN2<OFr^@S_<ab:6e@>e=7wF�~=j�8� 6$JU1b@gA�*ُ(�,�:NhQ�`N_N 1\�`&Sb//f��K�,N!�N#��<w:N+�N$O3�f.	g(u$
N"-N#4Y*\2�_5�m+1�2̑��7�4K�%O*/f g7�� $)*N1�N5bpb3Qe5eg05u�v!�,�6b�5�(�.�vb?e�l[ro�Q�v�&b�~)��&S�`#�b���� 7�N.`O�[-�_9bUhOop7zz<�3B�B�,� ُ-OOeQ&ɋ&D��:bxd_HQ$0R `S*b"�l%�3p���-T�  �(`'}p���p�Ǐ�N
�O��NN\#b�vw�#g"�v�&�`�b&	g b7��RQe }T0R�Q2�S"b"�eD�v(�9p���(�.�7�)i_	gO%c�pIQw��v\�$0R�v� �v�cCg�{)�_���v,{�N �f�%6R b'P��*�O�Q�v!��w���$�v�$Zb��v���Nc	$ 0R�b"Yu�v�#�S�v�$�*N-(W!A\+_ �_'b(�v�~-��-�2ۏ+ޘ-�bQe8x�$�O`OyY2bYe�v
N8N)N>pN:�O0�Q1�R/�S.�S@�S>T1�T8(W.PW:6Z=�`.�b8�b?�b<�b@cA!cD�c<@gAeg):k.�k6�s;(u6�y=z7�~6b6��5���Eߍ+;�Cj�A�@^�R��)Y�#$ N,�N2�N3`O40R�`�v6�z2ُ+�sQ&N\&�