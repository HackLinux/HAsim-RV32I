՞�db/)�ښ��B֢�.؁�h�\M�H;�W�Y��2�̨��IeΚ��(���;_,��S��q�AiD�}�dK+��8���f�����R�ȝþ�2�Z�8��Ә.��[�_��L��>o�#�E>�m��7s^;�>�?��`g氭�������D�,��m��F��֨ϼ������R�cN�'���VE��S۶a�������^�4��v��������xc�G�\�9GD�OG���w ���w���+�[g��'���]�L��NG'�u��������1����Pg iD��(�2�����v�k���5w���Q@�,�����'�����9+�ω3��?�H�&�ԴQX2����4	I���/"��
��>��V��ou�U���u����]�#l�J�]��r���6Ob{�3$�%a�6�%���'u�QA���]آ2�%���&��Mh�zҍ��(��j*C^\#��h�y�Z�=�48|��i�7�<a�t�Ʌ�$1������7�$ ����g|vn~+!�-�M�놥��R_���a( �Y����w�O�n�}���N���SتD?��"5L�����s`bf�49����Z*laT��v��7*�k)���������ã� ����pq"pG��g�ΠC LZ����|�ة ��ƘDd��p�@G�R�F�]�;B2|�4�c�m�jZV$z斵c*쪸��rfO��T�*�.�0���qeL}Uɻ���=���bm�5òv�F��ٚ+�&ʥ�+�V�/3�� �n�#\R4:��������3�ع�w@�5@ԅ���`qB�I)�ˋ���K��LG'+�������E̴j�V�h3��y�K�Xv��n�p���x3����X�isV`�x�	^���̤�y��FMC��7���������y�;�=ۣ���f^k�"������N�U���Я������V��i
V��V�n�o�O`�{ʋ�3�!P�/���k"'�#Q�&���%�4�1�ƣm�7���xdt��U�kޫP]�|���ts���?
8ǒ;������H{ĳ�b�nE���?�����4��4y�[4]2���<�(���mĸ�p?:,{�k�s�c�B���x��`�d��W��Ԫ��ro�ǖ��~O�[nqz��V�$�!���Z��'�c� pFB�u��pĩ&?6���\_�u�v&�0+�������η����ت�"������z���9��j��J��h�1hNg���l�]�A�:˦��Β���.���ӛ_������k|��X�=t�[da�g�m�����J	b�"گ{�����fTC̳��r�9e{���ߞ1�{A�^��7�+lx������J��ŎT�J��-�"�=/��Ά��E�k�d�V��L����%�Y��k�\�����l[ZhN�v� �;��J�4:!a.t��T`S���1֖�. F�&@���/V�#�#�9E��;{j�|�&�w���2�RȕH2���ӏc*�8MGS�`���Ԧ�R�����9IS]ϖ��T+��A�aT^Su���$e��d#����T�.;n+�*��j:�ԕ\>K
5�a�kY��bþ"-���_ӝp��æN|���Ŗ��&}������_2�|���_������r�v�]LP?+�9VD^�Mj́*�L����(N��LD,���z�N��ƈ`����7��b���F{4���eJ��n���ʇ=s�yxygdy�Tl4�
]{�=����G��������L�kq�=p�\��5ӵ(�>&W��rhi#�����_�0e���ڲ0k���pmb<I�w ��G�#|P�+)j��t�zIj쫔P�hq=r��e�߁���4ی�?�Y��3A��I��p��t1�8���ĤS�AscF<��WoJ�3��q�U~5�̲�r��'7:��j��e��9��m�u�u��M�z1o��&�E�����Y��bQy�Y��Omd3��ր6 iVbh�|'��n�{���N�ZbwE�a�*��7��;~��J�!�پ�<s}�?�%�(���`mF�
jcL��~�ĝJ�ڌ�}�y���l�#"[�$d�Q�Eg(
�'̡J4�����[↺h�;�=�c��,A�]��ow;�2�`��5!���t�Ԡ=^�8�8��
h.jG
5-T�KӼ�y��,�\.X��:����n�t����V ��Ȑ޾�$�m�\%E�5J�*���R�/��(����;]��}D��!����%��`|`d#<z]�U�9cVO��L��ݵ�i�K��[R�S�������sSv6B�d����k4^:�ɻ����ˤ���8�a�NW$\7�{���MO���G�#�&�Q2ǟ `X;6j����|�W�
͏9��N�*~���	����NB��ލ�[�%�բOc���_sS�����R(2*ق�fG�	��5B)=�9�P)�*�U�D���[K���+t�������_�"P^�C^��BX��g*햦('��+$���Hy��R'���~�o.ym��3w���lL;���A1��-<.�&LU�\$�S��ӎ��=KC?��c��d�c��^W�J9,5��m���ExR��ɗ��I�2��:�ɣ���a��F��#ò{m&T>Uo�������x���[$j��	xA�m��k��N��̑��x�)�{�������[H�fv|�b�fD����%DF��kE,�����U�;ZT�E̜�O��ckg�J|d�]��=�G�]�1���ɂ��mӲ��H|�i�Z��Q/[d�>'���~�4yo9�(��/���CVsG���\� ���%\��E�R�;��T�Ȣ~�a�9W^��]�D���1�G�,K(�� �zDoI��0��2ZCIIy'�s��c�S��z�~��t�E���?�������RS�&�̯-����"�MC0!1�8ޮ�F��v/�3�lO�Έ#�Ϟ��	�c�Q�׎������-4�b�����csC�Ԡ��P�+0��3oW�Axsj=P��"��E� ����|�����0��k?J�
���v��F����P�2�z�OY:����������xA���k�Qcz���L�̈'й,t��Խ�U�{[�C�8�{He0��`7}�̲֛��>�K��;�C��朴n1�$��r� �/"�+Ә]�NQ�j�z�e:.�+�����������9�E��uJ_��,�Ř5|�
6�V�ό�eu���{G�:���)2��q�0F��|%r�#ꦤ�y����Q�Z��������R"N,�Y#��:n+���D9$y�5�knٱfp�� %(��v�u��iEݨp�1��|����~S� >	T?��Syb��;�@V���'������A����2�'9��]�->fq�zc���:!̹5ye/����b{�ԄACL�}���c��/�R�ci�{z�M�I��}3$��J�^ �̝!]�Y��_�O�jZx�=���U�6�ڤ��Oa%�������h�F���E��k:��TdM2g�����@=Y��<����u�0#�Խ���?&��0������UQVp���ֱ��О).܁W�N�#"��p�o�b�$3�D��OR���Lr�loК��V�7�2��c�q���,�e�o��H�=e�`����'�m
2'����0�GGn�|(N����|� �	r �)�+�Eۖ�6���s�D7��W8E��fI�=���G��g����y��'i���)��Å��C��[��Վ�~*�f��Fܣ��r�{i���Q_���Z��w����6�����TB�'M�C�gDS˷i�'���fF�2|]}�}�+~�FC���T,S6��^)t�8P��4i����4�$�:�w5ݍҍ{=�*��Am0鍠.���B-�''�����k����1��o��ԩ6�ɽ$��!w��xe��\&��ԁq��~�<��Q]��ߢ�>k0�le����$���Y�.��%�b���xJ���7�mL�,yU��xC�(m����3��}���3�<��c�* Xf�d,�����[L�3�4�-���x�?^�ꥣ<j�E5Ka��lwKR�������a��!+D���&���nI���|��}�(/�_�7�ʚ��_lߜ��C�IQ�&ɬ*�M���8��g�Rx�����6����Y`j��msK\���bSwY�{
ꠛ�Tǌ����މZv�V�׽p�b���l�tk�أc��~�@���Gp>��G0,I���wZݻ;���������{f���;y�\Ky�*��3�UK�D��M�S>�� /��e�;��Xn;��/�k8��wJ6ǚ�D�]�ϰښE!Ki	j��:I��6�x�aؽ�2�(���;t����w���^F������E�

W��8���a�A��:mN�����������6�g��җ��5���u}��dZ�U  ��������]����AQ4��}�%.:��1A����=�E[�d��Q�Ot��[|�A�U��S�$+��e+E�C9��i9��q�綂w�����ģB��1�b�1h�a�r)K��<1!��;:����M���E��Tv|������F$f�4�B���|ޤz�BM.�N@m��L���d4}驡jF��Q;��a���݃���L����X?��g���"�4�ʊ�D��$He_s���ԺC&)��9�g�ި��%�m���^b|�sC�{�0JⱽZ^���Q��ӉS�Nq޼��'�f�|t��&�T�y;���"{��d��rv��b��@EpiH�U�{���t7u;3Ë�Ej����%A�v��X�c^9jYhգ�?ɡat�uZe��ܠ����|k��}H��M�T4��J�-� -֦A�=��M��M�#Ѭ��t( 6܆� ���2��_��a7���r��m�^��qj�ş�3��[���nx��|B�Z���#��jOm�x��v�2���В���������P:�JG$�2O��霅��a�lUۚa >>
��
�hֱ��КLE��7�b�`��iK���W�6f�v�>s��v���,ս�V�2��k�x�e�����ix��8���,|���BOM:��暣�Ý
8ʣڂr/�G��-�Hׇ_�U߶F�!WY�7��7�w�9�zqOc���MkJݛAZ��uI��_|��Cr���b�����\��~&��"Z˕���k�y��L"�fcsE^ac���U�-w~V(e^����;��f��oD�-�����srM�x�GȀ,7��i�r~�6&(x�,��:����Y-���l��tE`Cw�&78sV�0NG�<�b�nV�r`��r}n2{j�'-a
�K��*��ROya�Qل����^ϭ�Gz��ѝ�Wc��ǎ��X�,�����z��Z��;뤐~�Y�vVC�-���,�Yԗ�~x�lz��/�l~��uq����
��o���ȏ�wҠ���g����?���������l���\��{I���'���zd�a���+թ2��%��m9�b��
`�$���U'M.��F�� ��SH�T;�c%�ם[��D��"�����ɨ?:^�gEGj�BU���J�[%��q�o�&��_뫂�g��5|�u�G����o���#�=:O�����9�)�{����
����p����Ty7	�|*�:N��[�8��r>ҥn>�%/�Q�N��Oq�T�>�5Ŭը9��ˡ�8��m2\":�cuS+&��+��4
�"9�7^r�=��c�C�eb�ؤ~����Ks$�7O��&'�3�6�鞧`����󽢼�)N��MjM�_�<U~�����$�;B3��%��ͳ��.`xt�*��3�4��j���:ם��	�ZW­b��/QM�F�nc��|v���-&�3�d%�T��Ҝh�K(&/6QaA�H\l�.��]��B%7�f��r)1��T��'��'���4�!��wv�`vZ�ʲ�l�P��Yy>�i�7iuR2����X���{���[;�����A���".���"�z<�rV��ϔm?=���~����kq��&�	�ս��/�Mx��p����������S?6�I:/,_@������Tw��`���F,� ( `�ZK�4�V�SF4��}�B�2��`с��ߋ�!�ID�Ӏ"�n(�7�Y9�\�nt9�AV�y�1i�i@ n� c�m>s  H\��^ q(���` �*!�} q�~E�X9 � S�02��p=|26@�n9�U�{�}�{7A����P=zB�[5�[@�mc�n�a�w�n��2M��[�?��WJ� �z��6D%y�����4ExWU��g�v]yKpL�}��=B�4wx*yАL�K`p��GT�S�T���ѡ��
p�4 ��'酌�[0v�b��3���� ���
r���i?��1�!L�ܚ�_�J�lC���:5���I�/
^��`�y:��iJ���o�&�@���6
tD���@G\���z`��\
��B�|u��֛S9Pq� ����8��A"��j��+�_�P����kl�MtG
�*��䒯�(Б�RE+c�" ���DJX(Ԓ^�w�E�$G�Ê� S�!�&[G(�h�	r:���;b\�c��1D�� ��oK�Hcp	"V`O��X�;`ǈBl�O�yr�f��Hq�����J0#��-a�НF��r�e�3͈�f�^�-��a78��q.,NdT�-� ��pdd�,,�ង�f "j�B�pN�pKvH���x�p(��oHQ��*l��%ԑ�?�PK68��(���ѧ�� G��Bq8�@L�3J@����@�Č�K�3z=CA��*?�L��&0��ĬpD���IA$�A�?���{?LFLX���L�F�d����]7���nf疟O��a���`��&�-����l 6�h�W>�F��/0:!�����|�v����&��������\�sC�L����f?��(ϑ����x/7;{=e[�����	����/}�4%p� 8�ScsK�B���`���_��G�Q��[��/.�Q�xq����?�N���'�J��dɋ��%�q��'�����^@���Z����2�`�DT]DS�� �3�~���2;��=n�0�Fm�R�k��7 ϗ���)-y�m�p������!�{{��Ea�'�����C�U!~L���%��-Q�Q��`P�Q"#���<�{��F���.!��oC�5e�Y����V
����������5�n#���~�H)��J�ˑ���U�q���,�,���gب�S�;%ĦȪ]�,��r�4���������@�A�����u9�7u蘖�����5fgcȉ��k���B쁭á��������P�49_V�3-��{2�H��]>k�v����cO�鬗TŵL!�X�T�?�!3w&���q�L�;.����ğl�@��a�̴��Cmt'��#E�br,2�t���\�=kd��:|�t��9i��ל�]�eL�#��ZWd���ls`r�Af�+(ƒ�7O8�����<�T��]����!/��ȴ�݊�r_��*ͧ��$����+A:Ͷ�Cz���0������L<���ěV�.m{%�v��;�0%N������Z_�l {���q��r�畫;����#	�z�+�l�Ԃ���x۹
hx	�*���؍"*��'E�=�ᵳ�/;́�RY]����[�Ya΋^l4�#4j��g��peRDu"5�=�l�K:��d�x�GT�� >=b�U$r��p'��S�*C'i/uK��j�5����W�be�W8$[3�p���Ɵ��ލ��S��H��S�h��ͮ1tK`9A���+�w�XE�y�#��s�W��_��w��D�:��YG���Q3o@���$�:��k�-7Ve��g�y�Iʇ#��͵�8��n�;���Q���ɑ�H��C�j�oN%3���˪��w߃=��8w����ڲ����˯�쀗fڎojW#���שׁ���*OPz�{��L�s�A�����*I�on����Z���;�B�f����.����yu��¿�ͺ}5��7u�Ļ�\qǐ\�T�J�k�ɂ���w����)�?�\2�wp���V������6Tv��B�c���>a�B�J��[~FSZd�p*L�ld���X��F��l�+�҂�!�Ρ)��[�Bl(��8��i��c�
tk0?;����F�&oq�0F�*��nt�n��*����e@{��T�J��w���听�2���(���09�����$D��'��H>���?�"�����)��d���%q�g��P�_�<�)!q���|a
��'~�}$c��+X�)F����	S�%���|Sd��;�_��T�o��H��uTv����
c>C:��D�����z��I��P�(�Sf�GNՓ��u$Ǜ�[�C k[a9삀�!�Ҍ�<�'�� ���99� �iР�ּ�<F<"'��ut�L��EJ!HK��~=)�{��xm���01ٮA�ۙ���<]�L��-�0w�6��hla�7�6�������*\���>Hi����+��6E�6}�EK�ƌ8�˂�M���Ę�Zr�W�l���1>b�yT��yȻ)2�z�M�����V8��#XM�E��7o�ZF<n����j3 o��ൽF[x���&��`��}�H��,8l����"��[2�}��+�P��Q��S���'�&�^��C2JR�/&C�i�D����8��D���D��
�f��}?,�"�ʝ��=��]n\��C��O��Ŗ��sp B�8��;,��E�����Q���qb��k:����/�o�}V>��矾��,5�����&�~Jc�?����/�S}'��U�*�8������Z���7�����_�_���:���Z����Y?��t��=x�Q�9�� �����W��i�և��ՂkG?QWyw��C�U���K�k�?����W����������S����wPO���{;�����?�#�U���o�����zğ\�K�y�C�����C7Q9Q���Z4�/����'���Q�/t� ����x�	�eS�����^�YB|o*�&���!�T}#��^�ύ:�K�<%������kwt�����uh�@x/K�̈���ćJ����W��S ��oio^�G�;�?��|����������٦�q҈�|?r��U`f�J�ѷ������E�ke`_����p_�n���{}
HtXG��/��S"�����3Pg1�cE�_"�ou�'E�����j2��<��_�����:��)<Y��Q�crn�}<w�rB�����G���D��=s��?������϶�T���Ć�'������v��������Qx?�$�|�������`�4��Sݗ�s;�j�	�l$�w�H�t� ùu
D�(��t����}dQ��r� �s��i����7�/)�b��w:��g��P���������%#}{���V���Z�����8�W�.>'�B���S�����#T��y�̝�(n:D<�g �� y�Kw��l�,b>@#���nO��D��J.%B
_L��0�B���D�qM��ǥ��-A-�"��ˡG��b�UþzTi�^C��Tc7I����zR��<��8%��o��O8�s��Yޞ4E�8��G�q��j����l4O���}��U�ƚ��Ob�w�F���ƣ8|��.03?^��A�X�����^��F��C��1=��~�p��lm����䄺��	�Fk|�0@������t�f�##�)Yo��2�m�)��k-��2�.�׏��/��Nў"k7����l��xe���d*iRtl����^]���\t<���{�J�p�4q�C ںW�.�0ꦚ�f�%{C�B��]TBqe��p��}�V��c�����Ȋ12ٺ��V-�M���bRx�q���g�|���a��$O@~���.T�M�R>
e+�i���;MU
�P��!�r��yV���4S|B$ԗ��ؔ��.A�u��0�G����1�z�ȋ��V���>eW�p�Y��L��^����a�����J���7mx,pG-�`W2� 	y+��4�a�ro}u�9N�q|/cQ�7�����s>�o,;kt�Q�Ӑ۲V�X*^5//G9�-j^qWL�OQ^R��1�`6Ҁ	eQ��b��I���L�в�F6H�lX���I	�j��?��;���;��JҘ'Q�z Ӷ7f�n �c��[0�i�:��¤ҩ���/>}Cz�\c��ǜ��=F�\�d��.���q�{�M�	?WsA�1�H}�N�Ҷ��!��@��Hn�"d���9HtY�-��s+c��� %n���P�]EU^��Qo��L[,��P\�����{I2{q�v},5^-�H��F����(�i�]ŕ}X�<~�������E2�h�U��ϰ��mM����Y[k��y�� ]��p��0<�<﶐��S�J��Y�֘e詔���:w�`�nk��l����@O���N�qǧ�w��g�+�g�g������:���\��zB��4��*�&Tf� fU=��y4z��"sz=���yS�e~o5@�u����J��wG0�ʰ�������D}˸a���0�i;�b,�b�y.l�A����w( �O�T40$�>�Q/X\����f��Ys��D�I��ǘ��%��/�w-����d(����T�j\��P1�mY��7��O��@~�����������P�L�G�6\�L��F*~�;ʢ�����N�:\ykulI"~w��\99� M S
�� 7B	��25EpSD���BT>�E!2*�`$-`W���M��N{n��ڌ�<C�i��5�Gޞ�3��>��%�	��a��嚎Y���_:1��b�������F�)�8c�?���jO��3}����@1T�tǫT�
�)׹aG�v�Z��#wG_���b�mm�L���4>H����x� Q:�W���y�y�G��3�6[?E�|����Q�/Y�a�Z�Iv���|6�ݡh3e�I'�2}`r���<��ӷ$���}�8s�kLb���~�M����R�B�g��]�������@�w�oф�Gjȵd�
޺U�k���s�x
J�c��?�Q���
߇.�7r|O�$�_�?G�deR�d�J�d�R℘_tA,E�Y���V"�0*��"_h�Q���W�C�3�?��g����Z�)�|��u�����9��ģj�L�]	����b<���ѺX+�{��������G��>_:� �`L���F���62�65 !�_k������A�"�1���q��!�l>�6���0`��a���𵭦�X�+R�%�Y�S���~?N9A�K�����H��>���~o�?���{k������^3w)�����+��)c�f�#i��N柋x��W�e6vzY��φgz��s�Ĕ�#6;�4��vĴƂ���䗱}7��+��1$X�BWz��Ï�4t�c���8�HBѨmu�Ć�8ڣ�j(]OH `�x<�3�&���p����Tu��g=>�v<bq"=b�V��Z��U�F%CeV�Bb�4������J��bX42������d)ͧ�E�V�b�o1�����E|��|���XI��"6�`�F�C��_k]��4�`*�ݩ��;J&[zh�fg�E���7:�KMם	H9�N��ݪ�nl���fg��q��S<�w�vii�u7x � Wq��J���N��)U������h���`齁�(�gB���f�LYO_v���V�T�&7����U�h6g����	%v��
.���פ���*���˃a;�̰}�̔ᓆ�~�'^c����Lۼ)����3��@�G>
����8>d
6O6f:����	���TR٪������������U�V�c�G�|��jx�]�Y.U���$�
ݳg���{�k��x�	�3�խ�u�f���2z��/�D���^B�ކX��`<�n���̜�6����M6���lE�f����h�^>��.���������o�8����)�c(t����7�=��r����TtZHd�+>�����3m���b;=��}mmX��#�A���ט[J�9��J��߾\w �v�������u�_2����u�Gl�F�����oQ��Q�~KӣG�wS��ZI=��ޣ+r�1��v�=0���������2�e�z>2�� 8+L7�*�q�(5܅��kL+�Y�Z?���yљ�f��C��6^C&�+C��"�LS�}2���8rn�ܫU�^���ٗ�-�;��l�"��i���s�M!jy�X)�$Vp�W��t0�U��X���Q24��1X�H�������f8mL�����󙇾���T2�n�	��i(?8���r��]�&P?��_�6�`������ؕ������oH5�e嘖{pv�$V���w��.2W	�%��Dc�uoa���fQ��(��"���+In�t5fŷ�g����Nw�YY���p<c�[W��,�^_��t^6��u�*~�9E�������sK	��"غٙ�/������7��+��EH��0�{:y�f�xη��f���Gԇ9Z>P]Z�7�,K�I�i��J�"��֡�t�˝*��`_~�[��>ngٲZ�qJ�^z.�E?~�GI��.�4`���s��̹^WJ���C	\{�^B|�r
��>7zo�\�B⥝f]�}>1����b�z����b��>4Eo�{��3����}~�a�jEX��,E����E����%��*�T��6�^�ey��y�T��!��9�P�e���A���%+��8�7�O3��(�Ee7.?kZ�^ ���\p�M���E
����n�	�n���� 䣮 �@�融#6`` 0wO���AM�N�̠	�>�^n3%;��³�nz�=�4�kަȘ��=˵)~� ��qsU;��^@��@V��_��^�9�$8k��d ݪ�n����e'1�[z�D��Em�:���\_\�p��]�}�u�X��b=�f ����q�����D)��'��L�����r�S�V <_Z���C`yc�)�5e�d�&ˏ��p�*������Hg^X��G�&���#K#?�O���뗗�?��c9f8u�O�Ȟ�~�C�"�B��x���'��fv���A�4�om� � V2?����`�?�푀��8��a��J
-^a��x�W���߆?�S����-<���~&���j�p͜��E��N�U���ό���pmp�vokq=���L��b�<�SH�	ue�ݰ���3�P�G&K| t9a��y疀t�{Թ��oN�Ǻv[p���\�@�����N�m�<��'7��{:8�i��#�;��i���V�{�7����U�e_mȥ��җ�G�ʔ̭�D/���f����ݭ�|����b�����e�����k)�i�����f��E�Z��R=@�{,�*��~'Sޒ[^[EQ����G"Su��O��5��,D��iy_~�m�=ul��$��0H;��0�)C���E'�^ O.�`��r2��!Q�o�㥇�ǚ�s�ǽ�=�&��,_A�i�sS<kBk�,���Ъ"� ��I��UD���e��*�� K0É��ƪx��:�BC�:�����|&�(L���� zw�mGq4Fا2>�W�n
�+�׀�9yـN36���T��Z>'�K_lG�F8��ݿjw�d�ъ<����u�JiK����e�~#BZ">�a;Q>�7�ox��(䟸��d��|(�p�ʥW6�d$,<��z7>E�Fi�wr� kʼJ:��&k�'[]���S8��q^s�V���X�r��I���Toը(0�I�6�ߐH��o�HE3�%�W�KQ!d� ��A^�`{�:����u������7>��䅜�;������9w7�ш�*@����X���=w�#�D>����ZBdؽL!;ݩ\yES��~��#h���s����e �2��E��Ok�\��D��W������9 w�����<?�m���_��,�U�kU#�~]���F�~l�	�#�`6Z�X��a�$�I:�^��n1f���.�WxU���ן_{�_�G8���.?�c�w|��򾜭],����]	���K�{Z�\AYK����3�Q�B7��z8�G�Y�ϼ�V�Fd����&٘��c!��}Xes_���kL��W�0*I��g��T��$T�o�e��b� 5]΅%�{��b�-m��l��y2i,]99�{�-�ۓ֋�.\l�Bc����=ml��q�ۄ���";��9��FP����k�҉}zvf�8��`�u�y�1�����p
 ���@� �=@�Af� ��j`����f� 8��� ����Z��0@h�"3��!���r2�-�<z�ǝ�߱]��	���:P����AC���h�S��m�) ��4qi��q$�tL�7�'1bJ��f�JS�:[�U艢��$ø�ƹW5��Y�=�Xθ�[��p�!���T��_8�ú�ꓢ���s��ݠ��V~�8�}��~�ou�Y G�ŕ�q?Y~��(��	V;9�]xB^Ҡ[*<��g<�D�H�3&��O���g�oD�.l���|D�9�}������������QNf�����o���A��o8��go"�43��s579�:t:� @5��} �� ]�t�<���.<7������T!�c�k��wm���&r:���4�<�m��L�i�u��Q���nP��^�Y�f&Hb:�J�����������%]�3p�W�ѽk]^�3c
�{��mӜ�����f
�ׅt��d��s��?n��yy4y�"]i��~���W|;A(Z wd���K��,��H�:��.��y��5c>v�Y?��7c:r<��]ݽ)�<Y_��K)o�"'�]1�j��ǎ�K<���M�rD3�J�y���s�TL���FR����s�0X��e!.���Rµ҆���k\ژ$� �)�b6��N��tR�M[��wL*���y�%�gѕ��v��S��)���2�0pSm�ܓaW��Q�A�cK��U�JJ�I���;��q���qJ[�AR��ޣSt`���y�wK��W���n�$��G�`&���gn����6����ȫW��Y���֝��v�1��ջ��(2ֶ���I�!O3P���̆�;İi��T[���YU�]�y]ɓ�	g��},�.��]b�}�3�M���if�q�RkO<�^����(�EՄ�$�À�r��K��Q�P�Q�ؓ���W�-�� �Q�X�Ƽ?	��A2�ػ���l�>���X�ڧL����e 	h�� �&�b^�[i��}�X=��dJ�}���I�5���Q^{%F��q񲡛�֎���0sdf\�(BP�����9�vAb��6��볺��w�W�Nv��f�ϒ��aJ9<�)�J�	m\m̐Mkqm�:�O���I$�Q�z8�xms������{���{�����a>�1��uǼ�¿�i^�e%B.�f;-�6a�sXU`$�(��kޓ"Y�@e���̪z[,5S�z�����9��ąȮ�l�������Q�Pط����������N}���Ql�rRW|�c	�y�Ю�V�P�@��Z�<�ݟ �I�{$�7ݚB��.�(�s!�L�C�KOvf��FpN�Q�!�Q�]lliw�P�]f	1���"eCW��\��9�� Y)e��U���r�g��Ec�v���K
��Ah��«tM�kmR\i���l��dA2r�sL���NS�������z��+-8Jw��Ȁ�G�8��>�2`��&/�w%Q{��X�*.�+�����5Ǟ�����hP��d�Y����I`����"��-�7`�B(�P��:��w��[n\��{��OE�u��<���?�ӕ,2p��G�e��"\���A���|N񙶚kz%�@5�c�O ��ؾ��o��������b�N��S��?�?�Y�aes"�n�
f��^�A�������g�A���H>�� �����Mp�g�j_~k�|���
��- PGWM�Y�n�&��8�j��C����7�?��6Vy5Ƙ��x$��]�K}-)�}�]���U��^�<�DEBQ���dZw���!ʄp�O��~�[��osg��c��@�A�^������V�qJQJ�lK��u���W��u��NH���i{8j����k;��y������F�.�k62Q�z��o#�a�L�^�>�I �< �o��7�[ ��w�8� �k�~��������^�W?�����<��	�'�<�!�����X����*��A?����ߋp�Ņ�<)?�/,@�e�M���+?��.�X�^�Y����+��E��_��*q�޶@��<�]Ѡm����]Q��s��lW��峽��ˍ��h��,d	�}����m��k���ȟ�7�/ �cK�sr �;����?����|�{W��EN��r�z��~�51�����s������|������o�t��� ���;D=R�c��hO��udx�3�d���D7ڡ4��{�r6�<��P4�e|��'%�a��;����f����Ѩ]*�!*�L�@="�~.����݃���|d��}�d�-VYS�s IZvG(nڒ�=�j`��v
Z�qK��E_���@7O��V���U�����
���`��[����F��(�_�߰��0��W��B�YK�=I����5kY\����EMG͠�K��դ��R�����w�����l�˗/m�=���E�(E%��P>��>(���!��AiotNմ��ckǽ���˔O؝�Q�z��,3ڽ���@�0��Ȩ��(5G[򝩲)LG���(����rWS��f�sG�G��<�G��M�9㬅;����P�8�y�emo�)�h�Z�{�ܛ��|0��pMm�T����+л-�G���["�_>�|H�ԫq�&����p%�+�㋜��4r;���&��Q[��D�To���aEX��G�]�Yi�d�a1��^�4�X4) [8]��Q��S�YZ�P~� ��]�<$�q�t>�Za>���ɡ1c{���Rxo�hk8�a����>c�!�֪e�"�搷f��;-�"��٤;Y=�my�Ee��c��TU	���g�tV����4�O���>��Z���Y��6�ݼB�����m���u��O�����N��c��np,<��_���)�[���zD�c=?�3K:Z���]�,�wr&_׾-�R�由������K�������=ǪF&�����x�.TO>y��
(\�\?��%�w���p�+�*�
���V�VA,�÷�˂�"�=��(T�2
H3��bD ���
�J(�ug��l.�fb�GGt'�-Ve��l���DI9���8�2A�X�W%��J��)�U(�p�,#𢾇�d�6���H
R����-C�'��J�3ϖ?�`�����qj�#f��q=Z��߼fc���=�Y_����b�qX�"���$���a1q8,&�Ŕ㰘�8,�-��,�8,���8����eq���<��2�8\f��,�jÅ�b$p��:1���v�?o�I
�0<�4H�pR<\��
R<�L�����["��Z�ž�R��?1`�����W_�-q�d��4�p7�6������8!h���L8@F���6�	v��H�a�)�-�[k�۞�mO������ �Ɂl=s.� �6t�L�M&+������L��N������ w��Ͽ�}�{x����^����o7I�鿤�r�N?��Vt&����L���PS�Yr��cq�{����F�>9_��`^KC�?3_�k�ڄ-��!�W�A]��r�}~&K��dU57�d[k(��ء�������"��BT��ճ�pWF��!�&e�耍�������~�9��؜}%����͒ �'Umd�>'���}���QD����ke2|��%�qc>��F��o���M?�O�5�Y�>1�R�vر�ܕ��ne'UՆ�{ne~Q�Ї��[����8�B&���]A�Aan��w�K
�n5ݴF�p�<=��?n2��18l|z��N����\J��
���)�O\4t
�(J�f�i~�g�"l,�%El*��������Գ�Bf��|��$Ou�kF�}�'t��.��VC\��Ȍ���M	���I�<f��O�=R�dm���V��w����N�2�5��Q��Si�C>��uԵ�в���Z)�V�Hy��Օy��e��j�V��?2����c|d*��Й��q�Ⱦ�3(��ѹLo�GkU?Jbؕ���vN~1�P�z*�žzUpmx%jRXj��f��0��"U��5S9;�	�%X�Z���ʥV6p�%�ݩZ��3�.�HiK|�w��~Ȼ�����tmC^ޝ��IE��x0(ߵw����5u%�sǎ��"����<{���αIټ�$��+�ԛN��|�Ĳ��SdO��w�Q��t�̪Ǡh������&u����m>uV��=ɇ�3�#��C�({S��Zhk=��,\�:4Zn��[{�S��Xk�_d�d�!%���&vH��+�rä�k�̠�JX�v�:���D���"jt���*�$CS�ЕP�SuQ��QԸ=�%R����xX��V��?�2Q5��<�G&�;��B,1x��ی?4#�M���S�U��f�<h府�����>����]J���I���w�f
ٙD�����xx�G�ͣ��K��i~K|��7�jh����5�W�\} �o�J���}:�OSm&�v��.x��9��4c�y�m���C���!)�@�$m�h�!ȫ������Z���Bg�x��ٳ���!6�1Z:��o?J�ů/�M�evb7OZ2R@�Ϊ�-�",Y��GP]07>�t�f�G%qd�Q����(�=��r��N^��Tn�S���3!9'm[M������}�pU����q�Ox� =��S!��*��r����!�3�*���O<[�s��2��ܹJո5X��Sy����h�P�Z�LH����{Pg={P������I�<=^P�ʹ$�;-4c3��P(-J
���q̠�WTgH��bs4�����Y/��I[_�tn��޶ޮ�6�ΣP�BO����)�{�\�bS߅�G#��h�Zn^%��1mƬ9f5��(̑��ט3>2�@��uUx�����\��T�jh\���K2F(3�����n�^��.�ّ�kL�*".R�R0� 9ˌ�ծK�68V�^���	�A�/��Ͱ1 hh4�4<*H��a@�nL�������y�����cъO9�/6��ޑ/9�a��F2�c�4R���n9ІIj-t�k�H���+6A8']O�Y��i@�;3薏'�ګ�g"��
W5Jܥz4׹P�.C41�KsFMT?-~E)9�xܘ��r�sk�hl�Y��yDd�I;,Wo/ɛ���.�[t׋L칷��eE��P?:�5�K�Ж]�l�U}f�l� �Y��#�����Mr���[�/�9tz�����!.V
a�#����e�&ջ��Y�
���Ӌ�0��no-t2�Pk�1:�?��Dr�Q<zI�ۥJ�hìkp�`�l��yla�&,у�	�@s���� ���ݐ�t�m���tq�%��rж�I!y�͵g��G:���:�P/.侸_��k���;����n�ἐ]�%"�-���A#�X���uˬs�vN�mA3��]s�v�Iۀ/�:|}d�֞G1W��L��J+��BP�A"�27ьP�s�b�%�4W��IUL�b$_�T���]K:>XI#�ގ\E�]%���	m�I��9�X�~:X{�%7o]���l��x.����赱�d�&0l�*$*����:��,6_����Ks!���H1_���@�Ԉ�*8k��@N���!EO���?O/��`������jɟ+"ϼ�Ҫ�F�E)�5V� ĉ��~8��xu&R ��α���	ȱ�	��d+h�D>k4�J·��~ħθ��h�F(ں8!�gm�HGkQك�k3�'�����Z�7�ˊ�罋k��OG�"���_ϓ��e3O��Z�ʠ:�f������ ��,��;��%����{p��ww��{盪;S5u��;?֏սkuUw�ګ�?�������G���pq���g���x��sur2�w�7��燰�?z����/mQ+73I'#;�	�Ota����_C:�k�f�������y�����-�?����j?��
��?��k�Ӳ��S���5�}m����c+b��@�Z?����JЧO`x��s_]U�p��<�,>����h�W	1����~���z��ȉ1�z���a6J�j�f���v�j|:�d�y�ɪ�w˥1fF���,���G���M0����}��?�}������c��e�c�{�j������"�����Q��I��%y.;�E�Əޤ{��eNz:�� ���n����8�Ra2���4��*��4J�5�M):�!;�^A�bxwj	|��M��:�} �Z�J��q�� d@��s�y&�1�D�@���!Y��g��,(i+�H�\u,L�������bK�r�;��d���dy�@B��E��9ψ;058De�Xry ��@
���n~��n��TB��-���A�o�Tzd@�������Ri��&3���ȭ+u�N�R*�y��#�R����A�S���e���_��]���f�1}�3-��o�vQT�>s�m!�}��H�,�*�w��%��#��Ig#_#6~��7��d'�.��n��$�)�=B����6�T�u�I�I�c`�1�c�����ohWs�?�w��݉Ŧ;���w������1�{�\Spu�1x�/��tgJ���i�����'|����u�\Z�o�÷Q�i�����:�Z,���Q���~l�pz�+���;w�:�o:q{��R8N���g`��ȝ�>� ��K*���po�Ͱ�v��T�Sy�ɚ���n�[c����`R�h*�~e���'�J;M
{g������- o���	�ɚ�J;�W5b`�5�CsR�g�6u���������؉ݔl�9-�g�$��!�`N2�t�x��yfgǞMeΊ�f�݃6I&w���3N��y�ő�;[���g���,z)��9"sEd?��g�F�����Jcaò9�A��ʅ��>d��f���]r��M���N�"'��c�Jσ1��H��1�R�j�V���ѓt�%࢒�i�����}��5i�Ѷ�/�I�d"������l&�p;��U�EZ�`&QW?N���R�qsǈ!���|�4�N�|.p���{�����c����jhV��. Ֆ���O����E�-M�/M���3��kq.VV�����XX|&��S��V�@��=[��!���f�I���5�����>SH��Қo[A_J� ��1d$V_��A	����y�����j���o���t��,��1�rZC�����%9z�/��M}�o���I�y�kr���/�)���ʇR7EJ�T�hu)�nX�½�^��L۶'m��_ f�lm������덧����2��tVN~ E�{F�o:��5$yExI��2e��,�ԻPI��:J�.ْ��n�-d�j0H�x`�D4���"$��O,�}g��!��Q0�����Y�R3�ɘ[%}Բ �*rW�L>��tǐ��~�2N]��ݘ:�ݼ=��Kh�Ef
A��w$i�)yb������% �����X���R��9�+��+�ҦV��}���3.(�+(�15 a+:�|��}�)!_�9zk�$c@t���Pt�GY�)XX�mT��@�\l��y]m��W�%��E��^"�:��j�#X��S�r����YB�Z�\�F �k+�5H�y�Q�9Ά��-LF��a��Qϕ�5�ٜ�*&[?��s��F6K��w�W�*)�Z:>��4��D���O�zL0��ٽ����/��� *����j�R j
�հK�S|�?_M-����Wz'G%'��$��ۨ�~û�NO�f�>�:'�ɕL����+�8�_t~� Z83w�-��kt����t<<�R�;r�����&�{�%	�rl���� 
2�����T\]K�@/�Ns�����0�Ge{5e��v�r�I/A��h	�ϥe��������!��%������JE�L�|#�E[��B��4@��U���YA#�E�בО�"�h�EdE��⫝3�K�%7�ΊH��I����ֽ�y��6�o���Bl��T.��+�>��d�%T)�LA-��n�ϋ�3}��S�3ܓ]|&ɆS��8��I;�v=�Ϝ�����A�o�8�S�l�CE��C
sx��r*���=���k��a�f=����^�*cM����-�s%r�ϝ��7#Z���뾴%�����R��3�J��:����4��z���R2{p�X�;־n��q��C-���-���!9"��2n�4o�\K�N2�����64Nʢz��I�h=Q��8��Nft�	����X�	���'����>.K�4#�\�|C�G��B_�"\�s�W��\Es\B�K��0]�m�m%����=��W�VƎkַ�%�fle�G޾!౹�fw#_�"�+7?� #.�����I'[����N���d�S|/�KU��J��y�+��k,W�_\J�3�yR���B�����I�t=�Y��f�G�q`�[G����NÃ�aC�``��sz
��F}ͦ�c}(�s9j��$���v�L�#�0#���'�0JąG1���#�� ���7�>^.΢H�K�B�@�%DM(��go}i�ȊĸI�y�f�[��py�%p���k�f&�fvN�M>��7���Q��/o�Ue��s��o�Hwc�,淥Br2[�9FJS��Wn�)�/`(d���W�zkQ�9�a*8=Y�}�28@h/DBF�$�f��SF�U�%/�>$�7�o�"��+��3�
�h�Չ�"$��`(ٕ׏עG��<DXG�� ٸ޽�>* �<��nAk��]����'�؆�OW���H�������Ϡ_�s��3Q&�Ϟ7�½n�v�rw%��ՁyǙ�&L:�M�i\ 4�U�����N�E�{l ��Yؕm���J���ư�	�L�yєS?K�ʖ�s��o1��>�kH�'��(�A{�G�c�+EFci����8Vp����#8�_;6&UؖOp�����o�?s�p��[�~���DY��j@���S3�,�]k<
�U�l<u3��&)���y�k)}lqy�EO�)��y���}�	�x��%���RJ���ÔS?��Њχh��1I[vQ��e���AB��Y;�
C'a�,�-�d�شH
� f3xڦ��ᆲG��恟I�7�U�Yp�{��+N�iX5�q@���N�����T��m��S����Ӄ� ��6��2WJ/9^Q��'�����k�d��p�OĄo^k��_`��gXϨr�7VX��/��|������/�<�j2�x�����6��������`�Ŋ���/X�*SO���ZT�.��=6٫�E:��M��q6��_�B�q7R����|��.��74�q]l��3�B��P��݄��o�9�w��!�ۊ������Ϋ��>"��9R8�m?����GG���+l��T{D�"��=#�^�����=+X�ǨW$��qWŎ��5�`]RO�4�E��� ���AO��'�Ņmx7|E���b$_�b�{�ԩ	� ,�ϕO�C�K1#B�qK'}�y�F7��hFI��o�E
{��QRX�\`����ɖǇi���ȅ��T/p�xcv
E.u\�����2��)ݳ���ΚXۤ��x�$��y�@^g�x�Xl:���ɹ^(�y����9����������m���SG��D���iS'�����xI��Z巡�y��9ź��[w[�g\�����Q� ./Z孡b(n��g���8�S��S����
R.���ߠ-����C�R�'e짹ƫb��T�-����z���[���W��ۙ���zP�B>P�N������b�����e�G�A��,Hq�[mg�Y�;�o0"�1�PT��ic4�j��)��얮��|)��$�V�͒�w-�\�N�J�ʇ�U���a�r�+�Z?��-?3r�c�Z��"�Q$�p�/I+AA��O����e2���$��q�G���&-�ur٬⓵��m��#�n`���j�l�K4?{�}�i<��]lC\�^Q��M8�jYL��MvI2�i����{D��t���T��\4��ĩ��|'94~��G��Z�s�٣K���d���]����!��^LAr�n�b36�0�ׅ�����
 �#�$�KH!��f%�0վ�i�Z���@K�{r�H��}�ͷ8�Y���u�H�hؤ?"�i��l�3��`�m��KE��}h�r�K��Ҙ��Q�$>�b�K�1:�k[F�%N�iu�Gg`��
�5yA���I�����m�:��~��H�TӦ�Ͳ��a�G�΀f���GI>R�Z�Q�Y3���Ԑ�lZ��0q�O�l��g>C#w?\XϷ��/��-Xޟ_�V��5���A�z�
������	}Y�T����eF�Q�bX�LX�(D�����ȣ�w�c���*�����1$0�E�}z�br}&JG�e�v:�nVnC��[����yo	�"�	/�R��CƯ��MvB��P���W�!�gc�x��Zc}�CUv�xf���嫤LTs
��Xz�J&,vA����F���}|q[L:�u�ݔ�-2� ��pwY�+����4Ɍ���*�ǎ��G�����(0��.*�Ӗ�	�����5�W,cpm�/���/�ݨj�u�bp�Jq��k�jTv�;/%����߹0�����R��X-� ��aƿ�V�j��c����C`o�r�@Y�5r��'��JEr��M�#�D�(���3+1�"�A��J4�Լ@IXy��7��5
;pj&�j��ң��%z>��Y�˝M�]�m�&�6q��\K�*_���f��9�7��qp͐�ڡ�� C@����O�5�y ��Cz��ݟ�<�|Yɵ��9c������w���GXv�������
����m��_4I�����B5�,�ޕ��MM��˲Sҋ�*�<�n����|����O�ʥVdnS��n3K��I}�����i�j��l�y��|B���*��&����2�����<��#�F���ʮ�`�tK�)P`D��^٧�L�US	Cn1����q�e���G��%:b�����d�5��G���I� ��e�>�|I�9`ֽ��,�C�c�X� ���4	��Ib�(�$�2/�_�>�|�f�0�g�/{�5�s��r����D+e�T�@f#����u��eP�G+�/ڭ�櫭��]V���vGZS5L��A0ʄ�����X!(�m���-��8�WOk��3��Or��Tu]�6Ё7��x�[O�&#��G_�8�uy�s;@�|2t��9��8<�i�G|��b
a����0GV'[�(t�I.��Y�µ6nՠs� �,��'g��v�$�=�2�p.��"ݛ�z�j#H��\�J۱kbd ee�ql�;�LJ���������N�?v�c���o��z;���#a���8?ay�<�ɖ@ t����'�lh��/.X���`�f ��V�J���s$G�[�yz���h��}��t�*�؈#A�r��^��v�hn�
�94��5t�3�Vmn�a,H?f���]���;�����U��/��O�Qa`�y��\�󔸎If��� �/|�
�բ9�
�*rY�?��뺔���s����7y�6��6���VQ���n�Oސ��j��m������7I�	V^���Y#��e|�oX0�{8Թ�[ϱ�R:�$��`�䝏$��Yv�s����8�x��u_�5	��9<�.?ڻ���ޜLi���b����8,�!=�v�k}�z��eB�t����l�w1cЈܾ�WtB9�{wW��}p���[pp�x'�`�~�e�Pw(���Ñ�wb1����lB7A.�z��M4�FlמD���m��S�FaSr#[�-3hsyXaD���*���xm����6����1�;V�DN���cyّu~��J�T+̕M#Em�3�jp,o/�s�=��{�c7���Z{9���OGW�Ԓ?�	�{��&;�]�rqZO�C�Yf֝l;?.ɯdd�;'Rn94�~�OXn�a����e�g����2�Tgl)T����L������訡�r�{��(���?a}�a�^E7��bR�t٧U�PV�'���UV�'������9�@��� `�+^�ũi�Ŋ6�Ԉ�iEN�#��i�TJр�n�+pf��B,-�~n�4�&t�G?g@�[/|���ں
$e?��<�?/�u[lP�g�?�+�Ϝ��إ�5N�Or�A�j��w����E2�[~��ѝ��0�":���;�89M��$��5L�n';�����Kƃ�e�#`dr���������Y)S�j/�5��o/�?_�"���}�/�	]l1��*�bF�bF4/%c��'G�� �Z��F�����c
/!S���E�84/�8B���n���?_Y-ļ?O�7�bEo�����U2U#�j�$H�+DD:�8�:�2Ne��L��e�_���7l��۸\����s�^�=k"s��
���>"吾�2�0������9<y賗���a\:V���IRh�� �;�dMZ�d�Z*�����PY�z���H�7��y��Ȥ�zaNs��z�sw�'u�M�p�o�kظ�L1@Z��
�`��'Ǿ��oj�p6��T �i�[���^]0<?�V?ϊ_��6Uh,T�A#_�ˠ�
��<|J/��\��,���s��3�}�d	<� �9�h�=rG�j���>�x���SF�pf:cJ�3��U?���;O����w�株�Ty��a�����\���~�݅��i0J@A{��|��`�ް�Ԝ�u5��Z�cGŵ~'d��Y6/vm�Vc���vn�Pu#�-Uy��8��gאγ����6ý+���~"��.?3t�,�C�$����H��B��o�x��J�J�9�,�`���tl�2���\b�S:JD�=$@@��O��ʃƍ�l5�|�η�Y2lV�j.f�wj�;�'��fr�/^�i��H���{���
˵"�2!̓yz��\WVqK�I�ISMp�K��U7;rHZ�LY'��'�D�U��<p��Z)�n��3�;�{`�
 ��f��ٿȢ%��$�1ʕ�����v��:-�%��Ֆ8�$�)�>�=����w�L�3;sa���� \�A�{�ѻ��/���I��+78*�_2�!"sչ�M�^������Ē'=��F8�������(z�_���	���}��ʹ����`���Ҕq�<:��6sk�z� =^}��M�2x����\0 �B>��ՠ8arw/�����(���j���yb�g��X��ө�y�d��V�>���&�e{����(2�TJS��kK������V���U�������2+m�2��?��:���d�k��_��XMz���[��ю�%�u��u�a2r8�a�lC�b	颹&���e�VT���8�n�ģ��g�裵Z��%����qD���U����@���r�ct�jg'��a�H���j|�H=�x�!�jU��y*g��<f�:jM��`����7KJcpKr���|�n����˗&�)Yql�*����C�pb�Cy�?�qB��H�4!��N/��8XmO�ﶯ�	�M����ٞل�K��+Q��*�,�/�+u�yԱ�Q�Rs�2���g����N�a�<Do+��G�G��ŕˤ�񗪆M�l����\GN�s$\��H�9�	iO���=?��#t��s[n������/ͳ#'��n0���R3j�f���X����έ�07�?�mw�U!� K�,P���#�t؎�ƾR� %�q���4��;�?
�%ݯ�K���CMj��?�dH��2d7�?��↕��X�T�ڟ*��!��W��U����5#�c{�+�Z�{jL�� -u[��/�@V�j#�R��{��+����W��#ݸ:�ķ�@�����K:k����p$0�S��Q�h_zi�O�*�������o`"��W���<����((�n��0�	&�WHBF����A�0Vg'�@i�y~v2a2P#:_D��H��)/є�[x�w����G2�}t'\��?�M��k[*:�a$p20��%7�;��{��|��
w8�4^�./iI�u�!i�\��L�"���|�4�b��h��h��h��Rdx9��Lc���T���^m�L��|;��"h
="��?���Q�-_Gm�?4C����BY���RT�dbE,�R��{�;7�g'yɔ��p���X�E�☷��3n���6�pK�9�	X��9ה�Z��	�p�}q2������2��\��	$����x����]Jkq��|JеN�c��Km���r!Y���)\G�2�r\�<}8c8]�^��9���ibB� 
��3����:�O��H�[v�Q��>�!��t&t�\��H�/Bb��)z���S�	��DOWһ�����M�d��d;��?�ϐ�7�C!>���~ˎ��#���VĄBmq�'�>:P�:t聚+���~���/_������a������~*�ܳD��┤z�!J�g����rj�M��I �I�:;����f�P�"��#S.%E4�ņ�RR�"����Γ�ԓ�3阏ac���/2M�:��M���k �CK�uXV[�7z���-�Jw�t#Jw7��%]"]����H����t�ę����y޽��;�s]��w��k͹֜c�1��^����$y���=U2��dR��k��Y�
�d��.U���K�����'KzI��g��'�u�K�,�]��C�X�x:��m{~����}�EWY�$�&v�u��E-%��[�y�!�g���mnϺ�z�i*{qUK�t1�T��� ������_~�	�O�Pqv�ͯb�DG���h)X���t0�nD_�>dI���S8�=�͉Y��Vyd��ʷ��ڶ��|�b�#��D(�����E�M�,?ՙ�_��������j
imu�"�;O�[�����n��������ҧ�J�ol{���{x�k��LIhfR�K�/]���Yy��1ÒӲ�vxn�E�B3*s��F~2����\1�^�dZ�wtG��cF�T~��zYg+�U,�������=���.:���m�P#MC8��(*�mq������vV��a�6�{���N�:��u��P�"$�܏	�x4F�J�S#��Q�z$�!� 
B��'����nI�;\ 8����W���n�k�vb;6�0�c�w�ho�����	���O�ic�>ˑJF�I>���q��4�Q23��!^!!^�N���EXό�.�A'�o�W��:׬���G�&��Lj�p�z�u�ڞQ?�s��	*�w{K_��靕��N�{:�c��Y�-:]��Ll>���8|����_��d�a�벘�|�q,�i��D���J�"�6x��*����FY]���V�4Aߪ�G�� �#���[2�/�Z2�,����x�B4Y��OT���|o�>f��b��ü�`P�7�J[cބ+Io	�W��7�\�$��[�xf�x�?s�y�4�\6^7F����u≿��/t����ze*Uh^N^��E��)�K*qdp{�HF���"�S��I<�$/�[���C�,���92�H���P�x7�S�%���Ӫ`�*?��'��`���i�]b��u��Y�ze��'3��,���6['�b��r����� ����e�a�v(c^� � �;`qȦ+�Q�2��?o���0�J�ҩ�S/i`3�c3�U<z-���GX�1�ֲ05��ވ!������Hq��s���K�4��1�93��i/#І��S���H~ė,v�����ӛ,��^*��\N�gP@�B�:*-��ƪa��$3�䯇�'ߴ�$I���-?C<#��������Ȇ�@����������	ݕ��U�O_��!��w���]��b���j=��˟*~�6���;�YR� Y2B�
�Cp�$iM��A9NX�4f���ǿ ��q����a���,&��ڭ�!^!>p뗁��H̱�����
�C�6?J���~���'�}.�P&W��P���x�W��Lo�&����J*��'n�^`4�%AID�R��'�eu~��_�
�W���I��,]���<�+��)yw�0��Lqo#ǥ�#�[��~��eA����U��4�Y5��+�`Q���i��)���KxnR��4�_���VB1�b��G��R�ʢ˓�~��}蚉_���������Z�ԛ�X��!�ӡ�f� 5���#�a�i?TU�u����^>te~����6��GdîAdCbe������ų'���O\�Y�٧;���N̆'0�bg|��]sUY�a��,�m��3��=ʷA�o��Cm1.��Q����h�l����eI��˷yDo������X~^��VBG�+7�(�Kُ�r��r��6�-"7����2�`b����\D.�QiFh	�G�����b�3�xw$ڼ��LD_Q�k5�ܱ���YD4� ��K�A���,�9�<��(�Ž�!.�̐鯻�8���k_���N;��	`ۯ4�;����Gi�Ǩ����-��|d�3��8�v�;�ɲ&«g#���Iw)�则?�>;�ȝ�������T���˺�6 �	{����Q��]�6���}Ϲ�[	�i2!�8f�Η���yT�11�X~!�f|@ЮqDDl[p��n��.�.��Ԑb�֟�x�����)j����_�41���ʄ=!�|H�y��I\o�XW����7ħ2��h4�g�x�q>�m-3���}Vp�H�+Պ�k�:VS�������3��ߏ�~'���~PCc��}x`f��a����%�z�f=�R|[�z�C�����Uv�ٺ�u{����Y^fו���'f1�sG%��i=�(W�� 4q���/8��p�tw�nYMp��y�?� Y�`�� CxKF�S1Ѧ�i�gQ��-�o�p�Z����[y�0�c���H.���ZE�h��<t����������Ɛ҈�lָo�_}������
Gយ�ן��i�m
aX��\UEm��|��S��?�h�Ԝ��(@Ҫ^xq���gE��`�h�@����go�{���o/�ҷC\/��x��>m���`of^HrZ��$\Iv-��~{�/��/�(y�<��C���G�V�d��2��}c��v.�$�-^p̪N��2��Ui���w�����$|A�2s��;*4S�R{�~T��x�ߩ����La�q-��(�F�sA��n�k��#өU�����������U�>)�Wc�kw���vޔm�q��
�^@C�+Ӏf� W�әQ�qC޶q��6;��6��m����eF�gy�\��\u����o���f�Qp+���M��B�4uV����_��%Պ��܏&�$Y���Θ*��l��XB;�?b���V�+���"ytA���vB�����wɊ����lK�֑�$��G�#�sՊ�W���RR�F|��rA��O��N�u��rM������14mx��5M&�-ܖ�gJ�Y�H�?�ɲ��IdC��
7�^s��j�>�Q�v�Uк�6˧�R.��:�����r�reO�x�����0ң�c�N�>���/�K����vq�a�*&to���Ɂ�
H妢�B���Ul����$��5�a�Y/ەu���N?�ԫ��fd��W˩~�:�R���0&���zvD�o���HY�}������I���;F3\�ߏV#�QR�nTu�B \�|=�H_�Ic8
S^��v,(6T����e�)�����bY���J�>��wO���w��;�������@aV�M���56�c�$g���;��)������,�'i3D�Oك	�H���i�X'GX�..ӵ�|�Gc��$���90�e���zg�GI����6Z����ȾM��Y��=��t,CQ��y{�f`��{<�*z�q�U����:t�Ĝ����p��д�ރ��$w��g�?;�f�3��g|u|=�,j��!�Q�M�쫌hN	9Y=�����m>gY�3��_�^��=y��Z-��r�=\�Z���F9���b��1��R<f������#{��\�����gͅ���_��ۡ?�I�țڕ��̝���}j�|0�2�3�Y��QD�Ծ�9z(��ś/#��֦�+��bV�u`��d��k0�M��j�&􎷈��G-ߕ)�0��H�aL߭"%�;733!ht�7��"!x��Uu!c�x=�����cW��i����>�	���H!��0��iB�>y���=�p��K'|c�Q4�Φ���}����k=A^����
�����q�%Wl��ɯL"�n;�TI�K�/5�_�f��������ucD��m���9I���o���Ѹ�/d$/uEN�z5	�Nt�iN�KrZ!�H?]q���̸�5�9�z�"�m�d�O�7S<o����I�pld��^��e��J�8��6�aO�\;�~�f�jz�t7 G�U��Jgɂ�����5�����0�eJ���oQ����,�^�3}~n�;�΃>S:�,��4M����s˔�|���6�n��JxU;��׭^	A���_k����5�V��z��>��ԣ��?��,V�� 뭩����S��2��H��:�)�Zʄ�zu���y�O���+'QZ��P/l?נc����ux��m46�쥾Ȣ[�^�:��[,��G���&����p���}?y�i�}�~,�$M�ŮFY�C�n/���AE�'��W(�M�}�*���w��?��I�Nb%�,�.�	G�N�}��z��b���׻A�om���b?:��xD��|�r�X5a�����t��m��*?9��Ux�LHsz���qc	��	B����YךY�;͗���d��K���$uDn�T�BQ_�����<�|>���F����(������{�)̓��O8������;��-�_/^J��p�<e�4��������BVj�t��ueVͪ,؟���eɆ�lr!��G�N������m���?O�����v��M��[ڃ�8A���Ç�$�O���ʇZ�G�z~�80�P��!F<g�d~�FX���)�]|��-f�V���5�q�������Z�G�>;Q*�>����z��\��&��zS̈�%l谽�]��"۳x���d���b��Q�z�8VvBt�a?��:t@����������Xid,2�C��Tlp�(���g`����)z��[D�i��!�ѵ���B1v�U|���=H��q������3���U����u��Kсv]?���c�=}��u2QJ�\��P{���������򕕵\+���6���3���%#Q�����ޞ}G�5D����A�NV�Q��K<U*بG��*^���q���]�D�2�����6`�(l���QU`�X������4�:?6X9�M���q��izw�[����c���8}�_�,��&�-��7��'�p��G�v֍���ܾ���7y�J[�K�Ց�U�ЬW}���=���,���m������,����q.�����p�F)�t�9������������q�e���	>�s�:��Lc�ͯ
]H����.*1�,�푱�ÇK�n��5�������"�_O1�;}C�yZM��K �7��̵����&G�YK��~Zs��ia��k�7A:o�oi����yk�pA��r�����y��1�
��EX�Q������	pu|���bQ�~i��q2�b���nR]K��@��J<�-��v�#<�V%�Õ�]����7qV�z�l�����Z��Y\@�P��,F�d9O�dh��t�6I���ɻB��Oa
eQ���D^��R�v���I*6�mЕ�����ݛ��JJߕ�+��w�ɷ��Y��v�U+=Lsl��r^��ΐ��L�����S	:�8J��{V��}������ӟ·(?��T�D{J"e�\W,���]*?#�v��v6]J*�֏ǌe��i�d��&�\���j��z��,��%�-'�C�-�t�_�~<B�}�p�?�G��u}�7�s���ǙX���^N��lp��k&:�Y�_��v7�-�pZ0����W�G�b�a>7em�֢%��r�'#�˳�+r���MCZ�L�~�\�,)[tm%;�;6v�jX8�e����>��)y2v��?D���E���ֹI��iZ|���t����k��NK�W(�1��0C�.E)�)xߔ� |$�d���	MM�X��t�~銴{�����k=_Ed_�l�6V����������o����8�E�j��8�E�sHr�%s�X�E*Esڄ�EL-��ϣcͣ��ǈ*Q?����>òt������I�z�-����ǎ�_[;jH)ep��D���>9۲���6�����[�wQ�j��%�"��_Y��K�Iu)����Z^w���>Jy�����r����vW�5�]v�bJ+�pd̮jx�6!V8�6�*�C�!��d.e�x7F<��k/5.�jo�E��3�>���}YlXad��/��t�������)4I!���C�"ɯ���ґ/������J�s��U)Z쯫̂�>�V	q.���վ��6���3�D����\�����Z'Z7�Sk�]h�O�OH���%��ܯ�k.����bvp�l�6�ݥ���^+ j�8�ȧ"N��.��0Fbx�9�9'I�Ɔ�����t8�������Y&�kg8���`�.M/��`�7�c�1O��8�E�N)��N}r�w�)�r�[�����>ê�}��&rF#����EaY*Ol90b����|9F�r�b����Z�s����jC�����\���!qA�s��F����=��Rߏ���,�����G�S�2�(r�h^ex�?D����%�~�%�E��7f����ב�<�r�*�<�����5hG���ܝ�Yf�ׁ�^�p�S�����
��ٺ@�Zb������~�l�cZ�= �"}�-m�mVtY����� ��o��l��)���},�6G�U��wj��|�����L?�I���eS��t|R���&l�q�Kf�|n�RS�c�#ȡ��Y�g5���;)�)ZBk�P����(��7m�<�X׾!C+�3�!<��J0;6H-��B�K�y4�>�.'��{4��(��C��1e�Y��V�8V߽�+E�������s���,��K�w���YQ�\W*�aG��O�=J�)����P-��j?��������E�!<�_�ݖT�B�]�-v"�k��V��f
�3�y��t�V��~�δ�ݞ����ݐ��g���Z��|�g�H�FV_|�<nT)ex�@ǯ�<��:s�U�V����#/������YD+�����j�*7U���И��J��'l��XL*]�E�:�-H�9[��7�����.������zT�����H[�}�$�:|�^����H��C�2"vK�:{����;���R��:�̸>U��Q���D$}�M���Vt���ݎ�_}nF�ͽV3�议��\�iŒi�w���4[����Y�*�����)�"�ٷ���b7f��&>���#�B\�B�.��
����������9���Ǉ8s�f�~��=iU�3�`1���N��oVQ�����AN<��W?hv�2���^VY�R���6��R�|��g�����~*,��2��Ec�������F?ƥ�sr��fU*H�1��c@�}E��z)A)��v�v��~�oc�loc1��m�sD��pi��]��_'T���?7�W6;��œi������u[������ʬ��F�P�2���uK�%N��#�s ��]��+3s=:���Z럋*�,�ǋ��=��L`:�,�	`yޖ~y��q�+ܰ��Ρ����)�u��g�ѣ����q����lp�\«�T�Y�bԳ�Lq��/	W.�}�\�����^��c�RT����|[/S=�@�d������<B�v\�>W/�7V8<J��J�Y�RϦ�i����*�Y���Yu�{"83x9��8��ع1<XUʕGA*$��kx��Kz�r�xޱ��3%E�2�o՞u����*G������G�k���*��ʚ:B�SLє3���3���q�b��"�r���r�g����F�)�C�<��qO��E2ʛCA�����'G��.��//��7�*��I��v�^R�U���D����z���OКF����ԙ��J%���ZF����[V�M9R0�l�
����8@�D(����!�Y����3\���Y7YcA��%ǒ�h@4,ֱ�~N�~�hHXV⌜�JA�*��V������~�{��i,c�������p��9f���a�h�H��Hd��-	���yq�2���e������{��o���c�!��1��z_E?E�)�-PH�o�cҿ��󭃘�:%v7R:�gS��'-!��[�vTym�
b��c̏�g�.rL�����;�8�o<R4 ���A������<�>�	�Uf���ɸ�z���e�����
�j}���+�)&W�����p�E����ʦ�/~|�Q&��I`���ѵjGHX��p_��WVVԌ�wM$���?�k�%�;�E>{W�ޛ��QOX�PB3ӴM�ʺ#��a����L���������[�������?<޲�B�s�$e��!�V��0�YV5��c�7�H����M�3G�1	���<6��$Ү��Z=���E����r��0����́<��w���#B���S�q��>�u�[M�n�<ݿ�0Z{��`��[-׮��D ��6m���ϖm��"SYn_��)�#l%���w���Ubǩ�ǀ�ic^N{܀*S����W��O.�;�����J+	�eO�_dT�%
��u7.Z�Z>����h��*jt���a�M�oφ�/�끍߶��Cn%�eg�6�/+�dE9��cלg��B"�&/���by#��.����>�&���3z�=+h�,,�V$+bq3h,��w-R��Np�~��[n�˾yo�/>"�ӫlk��\��M�T%<B�����tV�t�Gsj��O������a>�0��{�b���}���C{O6������O���)Ǣ
����-%]c;松���~C
������JB=H3���'e$Q�}2�'4?�c��q'��s�_�N�>���;՘2��/��&Cr��}���,`�}��!�ɧ���>xj�����}�M`��\�5٘�w��
:q��a-���J�1ִ�v������!��q��4�u,���p)���1�ę�]b�V�;m��u}��T��4����g�N|���W�Z��<��F���6���b����d�c�C���=��b$,�#͠1����D�1����6�Ƌ(uZ����{�I��s�R�`.�,V��Iu�"�Oߥ[��<#.�F�=���j�<cNJ�R�u<~���/�x>�Lל�9�6|�:6���a���w���H߮��A�tQ����r�^!+J!R�`Ǧ����`@գ7��>�»�7 �gw�.ԝ���ն(q_V���ϙ���z6m&��{�u:���bn��\p/K+��a��rU��S�q�c�㒵7O�2��6Օi|[��|7X0K����U{�/j�2��3�|Z�b}��z7�(%Ȫ��}�rP݊��g���@�D�¨"�w?I��,Λ����f�&?͏<d9۞�i_CY�8�����S6F��G�.���_��n_'�;@���uC�Q�o:�����	��A�}�	Wǖ���̸�u!����tǡ� �'ʼ;*����fzjk,d?��y���ߴB�0�Cx$-:S�b1�Cl`v��0��ѐ�Q��p�r8�������`�娒����/��ٻ�u�X��'���\�6��#.�0|(M6��� �{2��X{ԋd�,{#*��pv!��j���bgAO0V�������+{*��ؽ�5�N4� ,�ywC��*��L"aAP�N�C�'���H؛��
o�~q&4��1'/�{x��=����P��C/J_�����
��{����|�1�sr6�}��֫P���g	��xk�٩/C_���u	^E���Bnn�'A���Ya��F��>"��3�wD�b�Μ��m��i1�$�k�hk=)3�9?�0L,�cr�$}c�wVb�KeXZ��k�;�;��y�-hx���/d�^C>J��
��P�D_���A�'���#6�^������x�G��:7Iw�|�ސW���45n%��pI���/��ڌ/O��
�t&�-��L�"j�?��yڰ~�!�?7�Q�!~rsJ�ĎLf#�\fcpQ����H�HF^����6�[m�O���YFׄ�+�=y��C��=���J�p�$Lat�}"�K{�}C{�u���渟;�qKmMq����Yw���.#�z�֋�&��q,�-�q���t��Q"�\&�k��,n��	����x�Iؑ';���+��戯x�2�WM������ L0�	?Yb��.�낛�,�Sʒ>�Q�k\�4������s_B�0dcO,����􃨘f��jG��u{i*j��{q�aa�$��-��3��7�H�*]�wI4�zW$�V��oH��$Z�ֶ��ߟJ���g+�_��I��)�{�.9h\�U�T��;aa����TXTN`�^���M�L��Xn�#wY�����dQO��x�ˬH�ݍ4��CL��d�lAm�ȁ�҂�P�����o���Q�2:��2	.#��9��ٽ9i����ށ5'��2*�y���1�"���2K�U���a�o�(SzN���#S��c�h��ek�R-���t�Fof���k����e-�67�����7Mї;�3�vEg�3L��Eߊ�vWս?Q��l
ܿ^�ߺD��w@�����M4'��f������-Yq����R�7��ХZ�����KU��gDNL�9��"4�Ke�-��WA�"|�q�E����[��!����n��G~F��c������,��坥��\�  ���ZROUk�b�1b�fg{sv�����qD�/I��I7���޹��a�ö��6C��T"���*'��7�� �����9�}�ݼ3 �S�K�n��G�~�
�k�������j�t,Lק,L��>�~��U�g�Z�������_��l]y8�t	��U����X�kW�>��Q��a�ӆr�A]����ͻ��G�4̽sX�|B�+g�Ò�Tz�*?��q�$�"[K���A醎�w���(?���{�����1�������T4Bv�➈�r��?��|s�,+�ڑ���I�蔃(�w��Bs̒rE��̓��ؔ�V�'rՏI�eߧ��z�E�?8���<�������_0;{����wT���W;!��".�e�
�g��RU|�m
ӜQ��}���ŵC>n����$���r�C=�SmՋ6M���2���^������zieo�:ɘ���H����ۻ<9�"м�u�����8zV�ܠ5��ǎ�Wǲd$��g��M���zI�tUyϝ�&K���_*�~*�sxoN�ew�唯�l��v~$�)�eY$=��������v�a�u����v�W$��KF�Ӡ����������r��K1'��x�Y����7���)ߟ��ޤ��9�?�_�k�m�d[�����Y�K�TR�	�Oo�@,:�L�����T�r��Z�ȗ��ȟ3j�$�s��*�i��u���1g��KK�ԫ��"�����3�T�Ok�#�C;�W+�������
�_�N�k�<ߙ��f�Y6��o]z�jv�GJY��8'8��S���T��T/;trϞkwu��:>����%۷N+��n��HX7}�"��"� ���������g2��+����!�e�<Xn{{���>�m�+�Xڇ{��;?�<���V���-)�vR^�a=��������%�����8�J�ȍ��e��u�����*��s/r����Z��y�-�p���kM�빝õ���Z씄�o�%�9�KC{_�5���o��pk�+�~��r�Tg��EmҗI�a"�����kv��>����/�Z��o3\Ky��q��9\�e���M:]�d� �Q�]�f�l�,1�*]>���cX�[�=o�k�:��m±_�K�*����{��ǥb�a�9��uo�_�a��%ʃ�X;���]���e|_�ٝ|9��:�E[=��ev鮹~��|>��4�|^�yc5�{��{����Ի�xu�e�uޝٖr�7p����N����0���l�x[�����v�>yR�'��&�)k�g�,�1�鯃��Ψ�͜��ٗ�Ӡ-�;\�ބ��]>�& �"��G�V�|y�y#���}��x=�)�D��s���8Os��+�z��y���\�	Uq��YSW�5[Nl��� �ƚH�y�T�=�s�T�ż���\�oL�⨖.y�����_e޸Ry��%b��$Ht�����݈.t ߸�dF���yu�Q��d���Y3ox�x��oH���׶��W�8Lu��Yȼ!ֵs�^�k=DrýYRZ�uq��lK:����+��*p�����4:�%�>;����5���a�5�r*j!m��n��&C�:s"�f�Ъx��
�I��i.٦7��c��O�G�J$~%a��L�;+����g|�8��v��C�|t-��O�a��00%�i��dғ&`0�pJ|�錳�{�����y��D|�Tu����=i?:A�D}^��Քe1�5��+1)zzt�P��DYޜ�А�:'97�#g��O�^FtF�"���dQZ&uæQ���1M��)<�G����i��Q�k�/�yL���{�M�k�>���1v&�"�a6���ѱ��,�� s#&�j����15)��s�2���|�JKK����]���A�C`S-�%9EG�S�〳������	g����+��X.;��5��]N?�V�j�=�@:�5�	I_|���n�_��\/<�UO1縏�$d0�j5.��fLMG���L�؛F���z��U�Td���=�o��r�U�Ɖ�&�������������Xƫ��k9z�����1*�S���C�[쏓Ҳ�$�|s���ӭ���S&R\�\�>Tڦ\]�L�����.o�|m=	��tYʘ��=J��_������i7?��0���k�)�G��������_|��E�6W�S+�f57<��:�?�<}�IU9e�H'�E��L0�R{�|WrA��=7��N�����~쎇����_Կ�;��Q��.�s��uF}�H5%L|���vs}u���ws�{w������v���^�h�Q�3��������=��
��椦�(Ǘ���!%���(��&E����W�Ka������fo-!��K�XVg�(���`ԫ��F/�w�m�6���6J��7,�_�A��D[A�bY1��|��y:G�K_?
����<�W<a�b:S4�F醑7��QP,�yz��%z���(�ZH\m�1Ԡ5d��24�6v5����*U���'d�U3�Bڒk/��>�Z�R�Lڼ�
� P�j&f �K���ɩ�p���
�f����=��~}!6�zx��/h���W0�s;���tծZ ��:��kVk@���OVB	<`�U�s9.���2ez�"���˹/I!���,��K�7� |��O��W���]	j'���{	�z��0|���������SFV���@�]跲��pÖ<���Zit���Sw����\�}�Am�S�kM=��#mn�������6w��R#�2�ͭ�@PH��M�2��ǡ2�dZ�Df��DXdN�`��$:ԅ���{� (U�܊5eb<���:\��b=g5p{��jV���7�T�:�"�n(�["x�2��=P]v/�a+�����	�_t���
��J:�uyH�܇����3��_ư�d�%�ĥ�l`�H3$���܂\����%�l_E&�&����$N�	������7�ָQcꄠ�bT�D(.[�*+Ѳ�j9��;K�ȇ_�@O��j~�Pt�4J�!��f������d-�C�� �8�Zl�G��Ro���	�4����I����A�1Bt	s�a�	s��k�����o�����\��a_���2�k �!}���5A�h����)P�"]����(1�D�kȜ�1聞 *�!ik�OuA�^ȿG:�ԃ��F)���Yw8M��-��E-kf�`�e�2K�~�B낕����
e���t��v��d�X�� i,��j%���=߃���G7�o4��������:���=��p<���-�
buދɄ�
�ܗR�f[�ƷbFȜ�q��,�\�����/v�i�dֺTH�ĨU�4L'�ʷ��vw��� s|�|Ex�
�Rѝ"Ô��v�ݫ
�_\�#�V}n�j?q	�oK�L✵9�@Bm��y)j����^��##�-����*-�,�m����[��v�H��/�-�I<W��\}��$Z����rK]�׉��BM��U�<�Y�\h�.:��m%�t,gZ�&��37�j°� .1_�����!����V̭�'[f�Q~T����{$ޑ�D��ԴxCQ�p���i�ߺ?��yFB�i���8S,���~�9��U~9d��p[7Z����+���~څ�g�K:�&�7{����%���^iR>�K�0�͔VuJ�Ļ�]�Wd�>�[/�6e�k�8Iz���#�t���@r��M�S�|�=�t��|��Hc�Hi��ܬ��{Ǖ�f���܏�O�+����s�;ʇ�����<�L ������	�ņ�
�`"��͓��܀��:rÂ5f ��ͳ
b,h����6�1,�,������b<���@��?a� ��5h�L �X{aA��`��
������Ӛo-�1�2��-���2Y�-SdݝK���=E��o���sƆ͍t�w�C��e��[~`u��&�\Wz�˷��~�Xw瘐[��e��[&��e��?�! 0i���z�pE��}}�X{�L:p˨ӷI 1��e��4�2�-�_�2V�-��2��PH��}��o��OX��-#��22�-�������"��P A���y3AlCI�e�ۜf(6Д��zPs�6�0Jڟ��7w<|ǥw\t�(�wuX0�P�{pP���*���Q(��� ���`�@�@9�m�6�?y� (�o��Q<�i��x��}Ar�e,�[Ƹc$����A��3$0 `����!F�t��䖱�n��o���,z�`M�@����ц��5on��1�o�]����9���A,� �a�_g С	���c)��FFO�c�^@���@���X� w��������3����2T����[FƾeԮ;�+G����#*�/�����Á�x��;�>`��C�U @���<�`.���s���٨0��2tǿ���O�]���=*4�t�~�O~c*Ԟ����O��C ��_�@c4�)E����5��� CP���AB��	�2:���e��[�>{C��[�i���[F�c8�[&��;�f��&��e�[&���'"	���;���;���[&s�e|h��g�������o����2��{�`��2B��y�-c���;f�eD�[�V��[���e����Nn?�	��2��];�)������� e�P�1[���������ݱ�-cB��!���~[�Ok&4n��&T~�����n��^X�q�C�O�\��8�i��;�cq��c�R,�O��2l������ ��-1�rۂqA����P� �cA�F�L����U��!�}�90
�y�C����P6� >�	:��m����@��+h��O V���q�����;^���[&{y�w,͹	B3�/@@L!ڻe8h�l�w�	�eX�;���7w\s�p$w�qˈ�Tv�XCw<z�8��Lx�:T�`.����'����;.�ex���1�@���	��Яo���"����l	��~���=t��c`M����*�^��ak��U����:ߡ�O��'�}X�: b
<t �DX��`�����s��灎�,�π��ψ�wx�>����6��׾�ȷ{m�%����]s��B���7�����n}{p�NA�����{`� ��Bxn���۽�8��..&��ŷwq:�o�����]\���۽"$�v�I���A���A�݃�����6%�őV��>��}�-��ܧ����(
v&F��/_�>��;lчЇrHFfJF6/��!�u�]�dJrl
Zlb

lfvv/�=l���5��^:;�54��)�iѿ��ޥ�^������i�)99���|q��I�Ws������<F��	E�����Gatk��;������q ��/�_�8B3��0r~i()�f�lc�W�� �+�[���!��&n��6�`��s��w����L���|�Y���	�}�Sp�Sp����U m  )�`|���_�}R�
V����+�+(�n5�����9�~.��n?��'����Yq�|�9Ѻ���k������g�T_���������t�,Z�ZgZ,�"��^�OX��p/n���������_���s��a)�������M�����̖�����]^C����)��@=���Zq��� �_�[=���V�`�	��a����_�Ьܷ�g�Vʡ�\�G�?���6��%ض��\�C���7w��k���|7������A�w�U�W���T?,U�_�\�7������I�����f�3�b�_-ȍ���?�����E�������ǿ�^��S���3��9��z��,,�'7���O�_~�/����� �����7��Sy[�˿u���?���?ן���������M�_��o>��8�/��5@��6�}A-	��U�C`�UdU��\��:����➹���!��^f�&^��c���`������`b�����to3<>і�:�Xu©Y����d.9��s��à� m���p�+E`��G���;�mW�-�sr3U8M�L��.����m��]�����	E����2X�~�w���pm�i�\�##6�y4Z����c��XA�lS����#'w����u��ܺO����szg'�Y��S��4�Nnҝ��N��Wo3%:,+±���0�2����I�~��N�qb[XJ�5,��z�z����khK���+�d'�P����w��fXȗ�4+z!��s�Y�vK�'c�Çf�1Z߷[W�)�b�R������;1��%���%7(����d���v����*�"�u	�c�� �)��Q���Yd�ǫ"&F� 5���/Bo�S���8WvW/���?(\����#R�L?��:��E曏���i,=E�ٹ�ߋ�sY ����n�N��8�m�<��~P�s?!A��Y*��!O���}���(�w�}œj�6?	i�Ք>o�N�_1m�x��D5���
癌��ÚJg����O�R<?�wUb��ޛ�T����&*q��븩��{�k���X%نnA��Ɏ�a+��iI�+���AIpsG*��Z�M�|K,)N�
�ع�>��߫�2�9����{lO/}L
O��tQ�;䧮�i� ��lCX�N��؏oI{y�s��y�bt��O6潲�$ܡ�C�����W)Y��0�YU�")��/��jg�T�< �x��7d-����֥��d~�ku �I�T�%]�#�F[@�4$�����|0LO�Q!G�[pw�<�O�������<�k��BN���y�C�7d�uCml��BS�rt��I>�Rr�ܴ0�G"$۱���u���K܄
��?ũ ;�M���#����0�5���й,y�w됙|�m=��؊��xY�������k�Z�|�Jp��_d�pu�'_�q�銌�/�V��=����|�r�����D(o�rW���=b��SN��f������V.���r�b'|$t��H�|���j���ױ�c�V���_I�gԭJjF��u;�ɉ�XY�[6�|�����nV��p:W���y"W���Ǌ�lpz;��Bh��Z�ɺ� ���t,��'1��|�? �O�5��g�$��2��r!"�l�&.��&���Vg��S�I�T��C�^����k���N��͂T{�(��v_4_�|�]~����?�h /�����Zn�g�;3�^d\�ZVG���7<�o8NB�Z*Q��������mhY/n%���r�V#�f=1��z��j�WY��e��{�>U8���9u�x���?��F�����PV�>�Yvj�u�u�y7�aY��Hr����%m���Ð�)jd�zߤ��y*���3YY��Q��V-��)���I��{K/�bT�g�_��Ƅ�O�v��.��cX��jY�S�-�X��Ak@%���W���z&�a&�+L�wA��i�[���R���*��̶��:t�g}�$����V�a5��T�W���+m�Ӊ�7]*.%J��QJҤ�Kۭt�é����K�����'LU��Ԧ\�� ��rH��� ��fG�WOV��-�x*yu�V��>W|0�(��5���ָh�T�C�#p.�ܜ�Ռy���EH'�Aǚ��f�Җ+`�Ek^MlQ=^�%�}Z�yu�*���������/�S$�X^��%����6��.����X���c��G����T�Ku��#Y�.v����~H�ʉ�;x2�JR��n�AY�Ҡ��CMg��S�g��Rў`�T�K�v�?��Y�t���?I^iI�7c��Z�q<n�����)�ت;����*������ĝۻ��&?�L4����`�=ڐ��!1�U��9���d^�2��[T�&�i���C�`���"3����<Lq��<�H�[���M�u�!:���׌�B$�Ci�K�j֏�6��F܊�S-u����T�w��~�������-�9W�i����\'�N`i�=��r?ae�M͏ςF)8��1�}O�Z��ҧ��8yo%%�j	?N��eݶ�*|�#tl+�on]Ԟ����<E5�SV�����R=-�2��ei�9�,�	;���y{�f�@�J��_I6?/d�lcc��)>�x@��jͳ�ȴ[wx���C֛5�Y">��M������y����D?�gP��6,<�e���Є��n�~M����}����J��M�J&���f�
�b��7���w�-iE��3-v�0��a{�p}��B�\�0fF�wO0
G�pl(�t�,��~�O
��]�C=�/9�;�1���(��롊���Ы@J~4Q��ύ<T([�£������*����Y��I��+�����??��U~qn�6���$�z�Cs�pE/*͒�Q�O=Nk�N%��O�|H�#
+��0��)^�n�5ih/8~�y�ɽ��˩���J��"�VߴS���^z��2�{�������s?=��m�#JD��r}�g2O���.���>һ�:��)�U�ʇkh���a����)鼔����SN�>$>ryM�ˋ�b$����6�U�t���n�\?x#���7߼�s�`���Å��gz¯C�:}��sȥ�.z��Гm���7W���EzH��^[�(�[�_�#U��,bVr�/R�u�����0Qt��տ�|������4�&�"z�ڭ��5N�QfD�~d�g��ki����&�H��q�6�����g�ÖU}����	/����}������I������P3YӔ�3Xdi�X.��"cPĒ3�18�$rE�I���6��mT��ʎ�:yu�
+�r���VE[B�qe��3�e�M���	��^/7�~^}){�x~t^�L��QR�L�i���t�GoN�}�L�K��s%�\�U�D��B�2u��x�y��3�5!ƣ�����Z���~��h�y�b<���hUZ��S�SCc����_䍹���|��j)+�2<
�+�5�͒�¹�����~����j��D���O���jV��l�0��2���^�a"�`817��/|��s���d�ںDe���(ک662)ۺZ}H{���WR[-�gG���<���:�C�"������ �����:�d�ϖ����.�5ͣh�u�k[�|rbQ3�H�u�.�07F�Q+�%��%��XQ�X�#5�����&=�K���$��fx��,�3���ϛ֒�\�>�7U=o�3Ԙo�a��z�w���~@�Υ��j��/�����i6��2ff�'�ҿ�(hd��75��M��g��n�n����2�C���_zu���^m�ӑH匰��$!�s{B�S�<JX�4sA���u�t�#gy���HSޯ��p�1�8xnb;�-�0%���:���[���[d/��z��k����I�/�ew`�ELp�1�����s���uͺuؙ��Y!"��R�*��uk��_�*K�ʾx��/rg�h.�U�8Z�i(2=��Bo�`�����Y<��0�1��02͟�������!y�`�f{�ՓY��UZ�o�W�!>����J�jDA���(u"K�֘G3�g�n-tH�l�4���>(�f����+',I����=��4a��Ǟ���������N�c�B��~��'G��r�����G�ʒRD�<p��r|͗Y迣^'J^�я$��~9YM����ke�*�e��W�O�H���/�)����7���g��&�W�p��[�EZA��7�o9L�6m<�y)��Ib�د�;�]��=\�v��G�.��A������XN��%��4�W�a9c�-'\/܏1t�}�"g�'��M
���ɍ;��]x䮯�_`�0�i��
w�v�n�3�]!��:=;b����uA�F9~��u����3�p��M/c�}W_��/�$�
��x��prS�]\�Q�����ܸa��}��B��C w�3:V	�k2#�k��K��fWZ�iJo��~xSX1`�r"K���> fK���	�"-)�w��4Da�l^�!fO$m�go�O��h�\�p��M�WBkt�a��e�战4��霨��~\�:W��y�a��M�c�b�[Z���ɔTF��z�o�6�$���4
�)�e��QSÎ�=y��(�>2��ě=N)!���
�Q�cs9ߏ��nG���đ����ĀX�"��O��4;N��I���$˟75"h����jTא��N2#�є@�[�Jo�xȏ�UQM
�T��
Q��1�x������Sҫ��ɍ�Ã�L�֙�1fӄ:)^%�P�j%z��g���N�L}/�x| ꎔ�L���u�&�v��9'U�(��\n����z����J$֧�|诌V�z�ȰW/��$�L�����]m�҅��~�P����`�@mV�n\Ga~��l��&}xyÕ4�����o�	�v��O-_�"�ˬk�}��7����I��K:���)[�ۥy�U	�u9�n#|��{��L�^G�:w�����}��"�|%�����:km�;�h�ܶ]x����E����'v�Rj�MlɱK^ì��QIS���<N�`�{�Y�r���G([úi���k����e�ye�e^i���?F��wG���ҳ��j�9�1$�,%g�
E>��M��&1�|��?��������D�w^n��d?�56����Y�)�i�{`��z��u!�< �I���=#X�)O*�;��Ԯ�W��^�{㜩��Yփ�:�V�E�Ⱥ����m"�.���)�f)���e$'B�Sˠ�"�ݷc�c�)ҝ��q���Lȡ��s�|<FЏc��d/4�g@��G	�.���]\af'��tK�	Qcb#7\�H6�L�o	�5D=���n=	ݯ�Qc^�:�(�/<@���z����>��PWӫԚӥ�z.}�ŰR��s7l��脌=9��D���O����7�4"�KyL['����v�R	4̹9����g�C��ӧ�z�2ikt~.�gE>�!�as;)Og��sS����s&xV:,}�V�A���Jǫ:BE�b�iC>C�z\a)a��+�Ka�����y�=�-O�e�n�&��`fç_i&�X����*�~�j��<����޿iqE%m���}���5��;��B��A!>bKd�zqv��W;H@��-;ff�����?)8��F+�k4�'��!+�2�9\��g����}��=U��5�h��DD���˭��ߊ�#a��{�Ym��ͯ��Hܥ1���(���,^���L'A�X+����W���+q�����?Mϛ�X?�/�1����ۇisi�<�n���@#�Y�xD����2Oi���I`�o=l��U��~A�s�J�F�5��2�u�����4���e���ݎ@���#�h�]	�I2\L6��j�	+X�I�Mu��r�]F�oV��<8߱VIRJ,)XYF-��R`�:��N�ɣp�^2���1%(�������U��)�	�8s�g[�r��ܱ�4Q�_�k���K����i��j2w$�l]%)ê\��ͦ�+��,-Ռ��k��/۫�@�����ɝ_};mw�D��-��U�ݘJN;/��ٝ��� �r�gsUm�K+����v�8��)���S�ށ~��ysΉ0����4��C���X/9�Ѿ�|�D�e�M��鏆����9x0"�t��잷�"�p�"�pQ��Y&
��6چ%���7e���q��#��uo�Xey��
�8���?7��Pσw�����wfk.��G8i��z��O�3j�7~e����~4�F�e�>��$��!���á4��E{S��p]�M^�'��<��`L�nĐe�E���8�#����t�g����i��-�#?0w)>	��g����\�*��/�h7t/o�7ek���:�%���B?T�j�'�b	�=<>9;��"Mp���ǡ�w����nn�qn�}�7m>C����
�O/:����>����D��b|��6�o�J��A��_m��-�_,'���=��)�;��j�<�~���N�����к�ɲh��2���为��ڮ�t�h���BB�L�1���q��P�� �Y�O���M��Mđ{���.�C4<68�b���m+��f�A����2F��$���ǽ=E�̄Y���g�?���Z��عx)p��UF���}Z�0J~���ܙ"/��Y�����r�z�:��L�s��y�d6�ȼ(�xV���<�Wt,�Е͆��i��#��U�hN�+CRhhx�����Z'���������h�Y.]rs��\9�Ĉ1��c�~���
�I�f�J|l;� �$E�%���YwQSg򩫰�q���4O���s;�+B>�$Xw��t}ٶ��B[8��9'�/Zӷ~�7U�M�-�<V
��e>r��Xje��e<nve�"� ��2�|������ߒe�o>7�޸b��$x�ȭ=�I���C�͓�W�!v����=D~7W����Ō��$^�~x�>��U=/��;Kڱ�T��S�6�=LW��G���HsO���^�:�o�$e�X��<-l琐$ixI�u�	A�ߙb�}H�_��F4���ME�O�Qs�R�����5A�(����Tg9��%��Z�[��JR6�W��2��7W&���_X@�%�fYK%�.��Ӆ�:Ŭ\��+�O,C�_��WA�z3������\ͨ��4��᎖`�I�[�AfRU������WX3�]ʟg�E���ӕY��֓��<u=�,�[\��_2�7��}� /��/�KT����j���-k�"���F5�T������R���(?PR�a呯�.����m<s8ҵ!��UӃ�y�F�9�bs���s��q�W�Z�����"�-�{	�i���>e��{Z��p:`;[D0#�җ�a��f�T)�h%���B�e��v�g��۶����lݢU6ݼZ[C�f�|3��mf�{-C��g���+�{y��	���W�k��&��b���!�w���_.���ކ���"���pN�t���k��4�ˋ����g�`�b�>I���c{0�=�z}�F�7�Z7OS�.�5�g݈���SLUv�6�+����Uf��L��6���DLfL�3G���4��hO����<�:�f��}:��u����*2a��̓��Ѭ4�'c��RD�x��3��*��0�H�dT#Q��]HѸS����{^SK�&'�=bQ������e��}�a:�Ŕ1K_�~e���2�Efm<�P���MvI�>��s9�_�:��OxI*�������:�<Z�53<G-��.���d�idG����5Tw�RΫ��1�*��ڱq���:ѰA�pS�EQ�Ew�AusAQl�s8��lY.�d�:7����ViL�"�~6�Ҧ��Iw��J8�
?��h�[5"�w��o�œ��;>�ظ�<�'���{�UۈG����(��+�S�sw��H_q�JU������M%�):�G��ʺj"ܤ�ׄA�'����p`��eӝ�i�r�Z(n�j�v������q��F̾��̓����g��i�;������_��xE����\�|H`�����U��V�����z�Tq}>��*�xr�0�=w�yZ��t@��
g���ޛ��8�������K��G�T�`V̈�>�D�"�0h�5�@W,�޺$���v�����ZM�	��׉�.U4�#L=�[6��/9��
����5�_�����,<{O)��~S�N�I_P����G��ա�|
�"�+�a�@�s��%��H�:^;�qv��̐ik&{qb�B�ϖӈ�K?s�K�`�K`���?��-p�^��Q.�������[�DZ��}W3�u�����`��oԖ�݉kKCT�&KeR|$����#�b������{�?~���[�����* �Nuʰ6��L��QaD����:��(e}|���NNCy!�'.4�
v�w������Q�f��4��M���;�y�L�O߿��Ee����!�5�yr��>�����3���3׏�H�"J"��V�%C=L_����+��|���@ֿ+)��������6'/�0� �*ǭ�~b���vC���J|�Y��D\��J�pt}_}�㵠��u���M�^ dt��%{���D����$^�qz+�K���]�SW���sl
�'AފaQ�D�;�>V���f�|x����8��-�Q�R����$^�>�8T��z����[�U�@�/�Fh�MXʽFY%�������q�G����Z���D��DO*)/���
_�|w�o<��N��������{Щqs.�_�>�5#�� ����,�@jIمH�3��EE��ך�I?!��� ���o������jL�H3�ol����L�_�Gzx�V�R^��\��{��8�� �u��3����"�7cx3	�옫T�g�aѲ��]��)��]5��${c�,�����o؋u���c}V�&]�Uv���h��X��Ž���TtO��L7w⎥��,�YU=�[.�;6��c�`�e%��m�1����R��i��dR��k���5Ƃ>�HZ�����F������h�y�+l�z����
�����(C����/&nh
y�]0�.���R��庤�Xr�	�	���6�|a��7�Z�>*����a�XȒ�E%���Uw��h���yj�Y�U�Q$5RE%}4�)�j������8MrL��?�h�ܷN��
���Ȓc��<���r�v��$n:'?P��~��5����ga�q���
��ѽ�Fqm���W<#�yo�z��q�T𞴐ڮv	I��ɜnKK�0�1�V8�|���"nL��[0ݘ���6z:��@����;���%�]�箟P̪�bM��[^U�S���n=:㰿Ea�Q�_�S� C|�3�pG�S^M��<۴�oȽ�s��"�K�E�W���oe��T~�_/p��Y^l�Q���/�拘����~d�m�I�E�������d�DC�rj>�B��b��e�^^���b�kÞ`��ֳ�h�V�o�"�	���#��L�?�d���#}7��J�K�hg��|-��֞�$9�F��ۙE�I�C��qU!&nŏ��@g���`����F��S�{�Wgە�M��'��m�L[l��ѻ,�9�
$^��[4�YR���<=�&���G	ҘPW7�6���h��P��V}�[2�li�z�,�����O�S��}1-��W�u��)?5�eq���.?]�r�t=Q������R��b��7�ь;��~�;y�г��Vw\�h<�^I�sAڐ�&ܝ�%�U������7�d�#��e3�݆����j2.�%��8�9��	ڤ��1D_�d�ُ��~d�2�Kd�x�a�q2��L�~?����F�3�������a��Y_��+��3bA^��]����5f�٪�����Q�!��a��ݡݑ�Q�!��a�ќ�����Q�!��a�х���dm��dn�}L�k	?�wJ�&i��gǝ�^�/'g�1dx|���zx�o�����B�"���Qd���d'�$��D *(���~\�8�<�LI����h
�^�1��I��N�|Q��mi5c�$���g������|3#9n���O�X`p@6�J��@���"�ݶ�cI��{[]�_�)���K�s~��-���5="m=�ۖ�	l ��J���~�*0Ma݋�j�N;]I*�S� i���U���]��H�+�6�C�9�S}�Z٬�Jd&=Vqrv�=ѓ�x���-J��E����m�ݕ����r�����ɓ���h���_k3C؏�_��Lz^����~i8���Z���m x��<ܻȧ�������}6���+�)��l����#5�T�W`c�� ��?i�#e�7nIz0I���$9��8}�fM���r���K�������
�q.�?�4��,�)����>7��B0���A� ���s���ܾ�����~��adngc������%�����A j�j�8-9%q-m��A��}�����s'���9������߻שi����)������)��������J*w�����Y%�%��E�^8�kh�IH����tt�}��.��?$$�:>�VѸ�YBE���\N���*i��u�����uĕ���ZFB��_�K�h�'i�i��	W,��r7�fp�qw<$yw���Ě���LCNC������l���*��wǜ�*�Rwǲ��w���)������r�w}���iP��֒����ri1�����s����ܾ���(���������]�+��{\���P.�^����_eFw:� �[��]򿕹ߕ��[�_�E���̿�kT�e�0^��(��{�1���̧�^f���e�:/s��e��{������C��?�������e^�06���K��e	��P��e��P�e�`�Dο����,�>��k����I�y�j�Ei`� LQ"��K; 8�(^���	zA0�ptr���DSg'gGz�������k40w�s�n#�^3ܟ���^V����_��d����Π�BC�!0����wA�ϻ ��]�������w���z�������8��@`�� �{a�/����[ D�
B�}�!��o�|x5�ѫ?I��,���
+���<RA��+�T"�M�W����vi�����T�X��D���X�b�m�<;,��A����{��Xy=���#�������b?4deYL�|�㕿�J����9�����_�����XX,l���m�?�Fx����`x��ѱ򘯨�%sޢ�
��������ֈP�v0�����i�����k#^t�=8%ũ�n�7���qf�EW���#���7nK�⢠-q��vbjRN%߉�^*$r��?݂�i�=�0��
_���mՕ�T.�~�}���d:Z�A �CK�}\I�o�9�$a"H%g�"Y␄!'�"ɀ��"YA%�I�* ��
HP� ����������[v�g�NuUu��>�οa��$繳��Q���������㟣c`���Y��*V��ڀ�\�Ri��b``[M}P���<<��<�^��V��jx{��Y��/�20�YJb���������>ڈ?cb ��D�;�&�$Q�����x>���4�I-�ʭ��+�|+y�]�m;�U����v��6�%<�D4k�*�ǒ/���>y��}.?���Qi�Sn��\�l�-]��-�\��:Z�A�h�Y;hdX��L�f�P�M�x�â9�=H�S�&�v��~3�i���4igVx_�d�� _�
ҹ�ǎ�MPw���P�4�z�^=}��0u7�'�`��B�	W6��$U0~:x?L�`I\�W��H���P'�'Z7��'�x���ֻ�*�5n��#��&��{�W�8=�	|f1}h��3�Fj�X��´�o�� �C&tN�j]4�o�"*} xYAԦHj�j�ԒP�m�yAI�CK���P)���ģ�Os�
���:�zq��)��Q�K���.�2�s,y/W��m��ORe����v:�9+��{����&z�x^�G2|�~��jӑ�Us_�|*��ٟpb��٨J�q����M��3=o0����������^��) m��������Œ7<����0�ǣ�$�D�g�w�! ��\�,nZ/���٤Ť2=z�(��8窙y!bcz8&=��:O��AP�-�O�Vf4�N(5�^ֽ��S�����Plx�j<�YI?U��p���1);�4�`������!�/e��B��.�6��:	q\����Rq#W���a���i�Q�:���3K��1�^���5w��7�n��<J]�6�?t�J�*`�{v���n�;�)��y5��O�
�	�g�����T��b�?�>q��y�떓�*��X^�?]��x�~w��	��-���=FuΊs�Cf"Jk�p�ٗ6_��_'��8�g�ݐ�����]�o�9[�[�w1����M}��/I�?ܯTɼ;s�y(2�������:j\�Z��{Yu����0�*Y�r�>�%��E|3^fIĦQ�y,Q����d�f枞,��w5�۰e��a����Gtf7<��"�V�s��aM0a�3�c'n����&l���3�|!�������"��Lܭ�����<��}o?�
��?`�3�|q��;�A2����VLQ��*���wr˓z��d�?5��9�N�jN� ��	L�K?ŪP�PK��l�Ŭ!�XƵ�`V2�0X�rFl�I�c�/�s>�'TH���p�K�a��C
;(o�/�S�M��Su٫'9%IMck>{�Ǥ�q�D���Kc`�@�y�O���o%d�Z��� �<C`?̐�`���ᐔ|����*��>�Z$�v�Á������)���F��  ��#�S�Z9r�i�-�� �u���?%���Z�k)����Pҟ��et&U(մ��-�R�#YP*��0��mSw���)�b�#L(�.�;WHz����Qo��_����E�#}>���EϜ��=BOj�5�)D�0%����j3��P�W�t���
4��Ma��7������8l��&�#��M���L[��|HE�{�27�G�"�r�_orT"TCt��K��O��d_C��/^�d��u��5��/.���{��0sS3�T4.�Դ�C��R��l[�Cx��٨�Ǭ��H����M���҆_�V�г�Z�ɯr�e_����|+�'?��'6X����:��D�~����6�\Wu��s�NQ#mTC���3�-W�Ιtthݰsڝ�f����]�3F:�	4�Ojɺ)��@����W�{T���;/�7�4����������(�WgGt����y�}S{�QL��1aÞk����f���(0D�ysa!��+v��bg,�8�K�33
s"j�,/U�UH{mf6�;{�Y��K�ވ�<N[��#�EF�-ݫ�M�o��c��l'�3��������Yd���x�r�G��/3O `"�_��D�Ք��/Lۧ��W	�ޏ�W7�u-i�%�I��s�Gڍ��f7.&�]ە����5E�m.�'�ϭ�']od9-.$v^�tT3 w�  w��˓�\��W��l��;�+!_�]%� ��5��.�����}�p_t��U8��*���W._�hN�P�<��[X_��Z�>u���l:^���O�G~��]ZJ����nZ}r0�p��O�ӛ�������F<#l��H H�#_�WP?���'�ȸF�瞛Cg�d��S�Rh�4i��З����������d8���A��-�D��/wK],�L1������*��<;A�:a��[qܸ��ݥ��	DEW�@�� 8���.Qdo@�ُh�F^*MZ<�9�f�}��m�V��lF���we��N"��8�^�@�n���]yW��)9�ӗ�.ū����}��p���}�f/�i���YF*dt.{����i���)�\��v�g]���rI�����+v����������*-����g�l���ϳ�-�j. �`]7��c�j�oN��o��W��h�(?�E��e~�W��7���:�K?��^�2\���b�"y\&z^���QvveRvY���:���]�D�,UH���6�hTC�ON��0��������e���gI���t*uZ�\�,ȧ�L������A�Y�Q�Y��Î.�,s�]��[����w���$J{O�]�9s���H�6DyBp�B��T�����l��H yZ����wIj_�~��F'����T��Ήtf����r����Ρ%���( �}��db"A�v�C�<)K�=���>�-R�4g���Khb{�
$�7�Q￞6�z������GK��^��w��Ү��v�'�=���e8.��k;h�pq�5�T������	U|R}���E�R��$�^ǥ���HMC�����~��Vgkk����_�8����&[wu���C(�\yoӋ,Px�[�P.j�v��_L�VW�:�~��� ���N\5q��*���3x1e�ͷǲuNr/F��ƪ�dQ��$<r���gx�ң� ����)Y��cL�Ʈ��������D�$)��^g��:6�����I2�4tZ0�$���m{�r��\�7��C�Zީ^]�Q�u,���"�s��L�-D¡����ד���W�������Oo�M�f��H��OyZ�x�s�g���U���T����v>z���ʋ	*l/�%�wwF<V��\ɘї��7(�~^eA{T���	�C�����]�\xBȜӥ���_քn�]m[}P����4��%`��i��0\ e�)f���z�d��A�k}�Y������j�@�P����H��MFY��� ��1F�ޖ�u��Xs\��U66�g�H�:�<�#8�+*g!�qH��8��	W5������O�w7dԊjM
�{3�����۩7ܞ�8<�m�G[d��e�x7/t�wU<חe���y�s�XsL��3%{&��^�3K��? �`�PCJ�d�]UUu�ưd��!�Ò��n��Q%	�,��Vt�&�
`���p��9�<�ڤtΨa�H)���������\�{�A��C��J��)M5ߞ�ӫrD�O
��/D|dŗ�Qs-b()�F����N��S��A�|��<��$��4�#|4�<r�V.:'.̇�}��pl��$6���"��x�f}ğfơ#���1����WR��`�Ȯk)Ϧ�H+H�iB_��ƴߏ�n���r
oC�66����Oyx�y�J��d�����!��(V���.+&�����S��Ԇ���يzrC����FW��m���2����syeOYCk��ש��#�=5�����?�X �����ߐ�;��6r�vm�U���ʣ T����%���$7�B��8����Be���&,����XB�\<T�SK�/�
�K��,���Px0�����"���E^�AH5i m�v��`�E˄Nd���!K��!��z�'4���n��V��A�Cы
��g��,=����1k����>�fa��.Jm��ɍ��1�)�Ϯ��u,&�'l�\���K�u7NI�-as��.Is��ڦ���K����'�K.M�u��e�rr�=��R�<������|p��#�}�ﮖ�f��,�v����r2�幔 /C�"W�75�r{�$z��^}��;(���c�{��sH�&���V����/�,H�<7Bj� -�I]�S��l4�B��	�<$<��9W��;Q��s��&�CLD�!
��ׅ��Ccѣ���Q�1�}�o���`�@��q��A:RHQXl�� = ��� Mb�^!�X�W�,�%��Z�Ŧo�|q&�b�ۀ�� H�`���xL ɂ��Ũ7	�ũ	�+�0�o ��k����]@BbpX��18��K ����x`Yk`�p����H� �b�{M@r���$��
�u� r~��F��A�i$>!H� q����G���8�(�N�u0�q.0
��DG������qv�0
3�!�,H*X��wLI�; (\��9h2���;���A�Xg<z0��)�u���$��!�����5 ��x�d�� 
���@$���C �"�CH�!������hۘ�Î�vǓ_a�S,���n,��b�~�pH'��{b�y��E����U�����a]�_��己�1������`��y`0~�0�x��+��K����`��sa0��e�غ�,>3Ǔ�p4&*|˯`�,/��
,���N���X�?B,v�&�,�/~6>�!X�^����K�G0��_1ؼx6l^4*xOl^M� a(s��+s�����ƂD�Ř����B�ƶe�b)�c�Q�s���ᐫذ*���,��c9�C�0�0m/��vˍ��8�Cu�|��a�ev/�����l7���0Alx ���Ŭ��X΋���^���^�/�0&�`��1b0z�X�`@�X�1�6��!�X~�_`8���cÑذ��-�&;
�"���E}��=����< #�G�4��S��&g�`��0�Q��X_e�/���a�|�Z�/0���E}'�!�_���%H�`������W�ѢB�����rf�C�Ժ�%��W��?j�C�j�C�Z�P��Z���O�mz,F�!��Q��P��~0�G�k����6t�#��Ϳ�U)G|�:�����xJjP<��)���3�$�K^���+��qvG�}l||��|6�����;r������%�PT�C��ɃG���j��3p< B�!@h($4l�3 >�
� �e0���C��� T)1xT�6��^�Q(�l���@�)C]"f��c����vb���~�o���C���Q�������,���� ���$�oa����?�W�������ǔ���9�ż�rl���Gc~�c���֯rt�v�튖���nv�LЎ�۾ɷ�qw�/�o��?��k��r�>;��K��*��?���l����灵�}�o�[�̏����[;��O�_��v�c[�;��_�Ͽ��
g������}��M@Z{_�+m0�q�cP��W���U�"%x�HO���5&��dWI"y��-b�ך�]Ί_z��J#�ͰG�M����Z�\.�����[��xs\�6������R�q }V�mK��媏+U+��S�į3t��Ρ���Q8A�6��j��!�h���w��hI���u��K�w
]���y�o��D&;�2;N0	�rVkV �q_3��;d���R��]���� xc� ��I��gz���Ϋ�fe@��"�y�	cK���ޛ�\Z�f�a��N�*/zXd��:��S���ˎǦ���,.\��=�z���*w��$)&���V�
�Y����_�i.4-�{EOH������ؖ�5�d���w�/�b~V%��A7';�m!��YM\	���S8ǭIx+�G1ߌ0������Ȧ�@��S�mMn|(G.�I-{�w�'@fl<^��&w7�x�Q+����o?P��Y��2�Qf���h�[��~�\u/j�K,W5��=�H��!���X�^I��r���s�<�]y����_�s��u�v �=�Y
gt���K~$����z�9孾))����&x��g���^ߎ�yqĦFVg��5����3��Շ2�'0�4��������b���5�ZC|����b�yX�A�Cݾc�䅤�n��fi{\|H?j���Kc�����B���?<]�p���k�+�#���_�^k���~Ǣ�����6he$�]�n���ϏG4�K�s�Z��T��-�	�se�}��Ld��k���_�%���b9%���O1y����4';�S����Ȯ���Uīg����4wã�����uS�S�����:���H�tݷ�ʪR�"ʼ�9���̍�_]�vA�.E��m�l�ŲJ�Ԩ(�ZJ8[������If����l��gW�y5���Vm��,�}��Ԁ�"�w�wN��l�g��[�%:�Y�.�����J��/�j�U��t��dd���|}X^s�G"Z�k������q��������$��p ��K��������*xW�7�9�������tQSNQ��1�ټ��fs/�am�������=��>8Ş�T�h=��7|H:g<DYrQ�Y\8���BH4Pa.�_�x8�K��m��P�Ww��/2��Mi�ڜS����>��*ҕP����C�x�v�:���PJ0_gD�eV�|���@e��H9�ؼM����$v�B4��N�����#�=�'H�yK�H����
%�v*��ih��ݬ���5�[�wL�퍩*�� ��(л�A�iʸ�P���,+����y�ʊ��!�K�ĕ
�7ʧ���$t~ق}LR��o�h=yO��!���Q����=xzΤ��q;�Fj:�^&ߔ��`.y��ͨ�-r��C]]������F�<�'���{�e�0��|m|}�BE��~_�]
�4/>]|�9�y�v�4,Α䉓%^�v4uF��P�I�:ɵ$kF�z�is���5ϣz��d	�Z_���r��7�g�$��OWk�	&�UQ���_
��1�MS�~��#+X�m6x:��N�!���Md$�Yʩc_���U�{Q������{Κ�g��ҙ�Lu܇>�*���?^�q@�y]yn�D������<؉{�=���GX�����(����
��yX�L�).�_��4�yҚNx�>_Z���譚���{NB�˾�Ⱥ��{N��+�	fZ]*��ş���Q�x�[א'\y��p�B_ĴE�v�=�����ng�k�&'˜�|�|�����I<��?�M��|�'awVb���W�C�<�_s���n�=��\���S�w�ަ�ʢ�R:ˑ��uV���� �=a������]-�������<�����(��^0�~�}I������`c*��KRd��.�'|&t텎�W���o�)L�0$���m=�(l�l�a\{�f��\�I�31�����E��	E�A�P�U�P��V5�5�i	�!C���O_W�W���Vѕ�5(����/|��ik���᮰��e�U�e�9TV����}�I����o����/�������f���9A��� �y��\�Ӓp1��m�v�׶m۶m۶m۶mۜp4�򼕵��+H���`LJ��&���:�Q��JH&DG�'��>q��G>��D�ݫeb>�dE�K��mLi���}i�����N͗����+�9��Q�I��K�I��6���":���	�!���`\��F��h
"Fr[��{�!��;�R��鮰+#˷�鷗W@]!��%ڋX
Z�tY%�vN>녪a$L����?��c�'�1}:���t�
���3Le� H�W�A���T��|���\��~���"h�	�[�J>����B����)2(�s��k�X^A��N�z�A�2��3���Fiu]�JoV��[,���ν��c�y����˛8U��Q�\aԷ0�.E=���E9���Z�҃
T� s]'u(�*�� �����{O �b�$�J��N�ܞǑ4Aq�#1�+W��{�1�����:\�+}��~�I�A�H5z�u�#=��Zuq�b2s��7k����n�bwDuqFR��@��~���g���Rf�>�Nnޢ^2�����
[s=��d{�ؼ CU[N�'(�/i}�&�.'jl��?7������l��/���I��+�c��cgC�F�_r>dc�;�`�r�<#Io���;�~hU��ם@�����M��%ž	*ߒuA��~t1Դ6�.�`=u�7N���k�f�s(������dƫ31>���HzŞjl4h9�V�co2+��(���t��/�33�n<uͤ��wI�\'���m���=鹄"v�o��Κ�Y�FY��P�����(��η� �Bj	�yߔ�EX:j�S2���˕ �(�[�h|S&�ݕ��%���D�9�/@�7�ӫ�5MC��<Ʋ^{�|ʷt=�bo�%��έ��:�Ғ���8�wk#<�L�"ꚃ饪[��n�Z��N1���bW��Ϩl5��O*�OC=zW>�POE|�d�DNG��,�d��z�>�	��ꞑ�\=6&�N����d��Z�f�HF��g��`3��g�!)z%[ɰ4�ڬҕ&Y�0:�L�ܪ}ܢ.�I�੝O����ѓ���u���ݧh`��cq�zԔ��US�3F.F��A�H��@)j�_r A����+�5��j+V�`pV>�����$67Nu���=�!��O�1ŗ���?�~\�R��a�����@2�'���Sp�����0|����������7�H� ��0���:f��G������;.��������8�O��NԴ~~^?�h�٣7���;���S��O�W����_�w����*oy��~�K�>=,m�������Å�၄١W��mO���]F���.�p�|��}�+��=?,б8s�8[�sE�gSm�k������k���:R��k�?��)�:��wؿ/8:H;���?3�~P��>J۽(#״�߳�"p5�ª�F�W��-+���X����յe�@}��ev_w�xo�
�!�>��$���g�ղsS����i�0y*p����$�>�x�%�TQ2����ijk�B��G��D��%�'+�GnD�a�!��ϫRa@08u�WF�pd�n=o�a%C������^5 }J��  �"C&�����#��A�l^2A����D�q&��R�sv��|�[�������n�����0��*�XJ��]1����܁��RB�W����H�_U�'��w'�����9�<��$CO '9eҺ�D��av2����G�O�,�m:<�d��)I4S(�,Ǌ������eb�Nպe�����'%U��?�;
�<�>�W������h� *��� Z��ƭ������Fo�8�  �}F$X~s'���U�ȧ�"#"��r�j1��N�O��Ue�s�����xnY秘��3,|��}gdg�]�v=|{*�Ye���k�EX��H�o~���$1S��<��lsW܌��qߨ�FS��HN��}�?�t��)�YK�~6#���,���ܝ5Ʋ��ۣӤ�M�g�{a9��<�G|Y_6@>�|,��ZE)"9$��
<hPWꂑ�Y�V����1.e/��1_�g�iI��V�	B�B���2ب&lXL�O�t��� n)Z�RQ62�����:�o�1��B�<��1�Κ����=S@{ZS�ɤ���y�!���� ���B����G�D��4�A7��K�t �
X�]3��w�}�'!�Egg��$	�D-�Hp`��.N��H����mFA�̜��NUZ9��o"_"0x�/��N�S;�!t!^4�! �o�������X0���W��diu��w�δ���ܧ��v3��K�756���ҳ��x��M�����1��Y��yY�
H~�z�	N��]W�W����7��ͧ�ʫ���$v�xt�g7��&�K;bW7V��S�	�}tž��:�O�7����������J������	m8��c��MwD^\�o�V���AO�
��7Ѿt3�CBn��t\�V�r8Y���e_�J���Ƅg�����{Po/I�p4�V�J!�ȸI�gC]'+�9e�6i������I
ڌ�d���P�o9�S��V�v>����䓎��fd�$Mߐ�A�T�ҞI�6��a-2->)������~d�$�I��N�v�U�y�̑���4*��O�0�}_�1�Ԇ����5��B��s|��(w4N��٫�S ��D9����c����ӧX��j�P+Ƃ�B�5�tk���DL����GR�_�S�����I�Jc9[���Gn}1���aZ0������<�6�� *�TlQ�������	���˯�ْu�x���U�5U�cL���{K�l��;���BWar�Yi��n�z�'<����
��.F^W�m���'��M:;��ձ@�!�}�����Y��%2�܀�X��k1O�e���N$u�?�[qW��#�Sǉ���-ȱG;�D���}Zi�+4 �6p�ֲ6�Õ����Bo5�à*����B"p8��S�B�c!+#���R|��{�&7-�-,���������'@Z�kP�w:�s�	\�$�b��C�C&������dZ�bV`TV����S|H| 3��v��/2f3���G֊��,ӛ@��c��[��/��_<ݮ�޺�+��6�ʅ|cj���\2/�~�>�v�o��1��ȵ����������� ����~��YbU/�Y����������[�pP ��N��;^V���	f��1�vc����f�c�z�=�rD=D}�?�|ڎ���1{�0)Sh�A�>\�L�7�+n�ӿ��}��׎76���(;���k�wp�%���T[��8o\��6d$�	a�.�o$m�2M.��cH�C�2�
�gl"���J����56�G�J�M���y����^�HٕV7VZ��\�)F<���K�uM[%�T�o�P7Q*�����	vW]�~cϼ�P����i���Z���x[5�+6���,2���k"�RE��V�8=$D��px�\1ʎ4Km��sBv��s�Z���ߍ��\����j3L��Y���>�����������=8�$�d��)A��i~�̩~��)B��g�0t
������5p�����ڶ�s��/���7����g�����v��� �o��X��j 1{ig�KI���`��\oۄnn7��m@��]߯��_���O��Hh���qI��u<���q��
h~'��lZ�)�7T���>��)�Nv�"Ɖ�s#������G	Wͯ��
���#Z7�vy<�����@�(��M[/��}fe|�	��ȆV{��v��'	@�O�Gu��6�G��S�������o�	2�[�:m�&�����N�'-7�j���@�W�n�@J�*�֕��Aܧy�S,:R�������C�y	!��Q�6Rr�P����M��Iu*�������n���	'�-*G��t'Z7�˦�%�Қ�ȵ��yUr|rt�غ�����e������wY�gvU3�O�Dx΂���il���e��(�{O���˿o�x�#��jn�fo����ͫ�����7�q�����& �.�=�b t�����23p�<�B���u1�������<_Y�b9n��$��a9iq����BS9�3�����5&KᎶ0�	���u�>�N���>cY��"�_?�F�Å��2d�C"����58a��H�Vbۃ�bO��Dd[���r�	nT�~�WgZ��qp�䗜XM�����l�G�������A|�������M�n+_߬Q0���x��0����kc���σ�QY����
ѷ�.��"X[P��u\��w��������es6���tx���w�ۂ�w�ϦO�w�xɞ��e~��"k��a����&��bL4<{��ɾD��+y�<�f���O�R_˴���oI�(|Fg�㆜�^� �%�g������X�N7y�_y:�����fU�����{!;�=�ԯ��c�UsJ�`�ZF~ˊ����(rr�j9�]��tǩ�ps[��U���e�1FF��GM��7W	9I9T��cq,7CW��8(��1��N�a���ɋ�@���[	�߉�����N�d���,�N�5�U~��ˬXᲱ�u	7O!C%����d�]��ϳ�[kbٺ������6�z��S߸�:�>G�sFh�X��.�i�}����۠<�䫼�x�ƽr���&���h�t�I������`�ų45��ܶ���{d	ۘwF���9�M�+D�	�u�J��(�$�Oܛ[��2�:��6�e�_eQ�A���7:.�@^�ϸ;�fƮQ���jGa��" UZvN���X�*k9�]{�����V�x.OQV�YN?I9N��{�Mm�	�N�?����Q��ՄhXc�Z�a�W�]xw�ů�t��,�3]�m�S\-���Y�ڄ�H���G�j�qS�ƅ�̵b}ޛ�'"r�@��5=M��(R4
�;N��5#��R.��YD.#C���OVm����Y����?�Ii/[�+��5��������&�Y$'����a�*�^��<u_7��Jv�̯�"0��p'�	��@��#`��?�׺;���ƿ�U��e-��dq��v"��k���������ƈ�k�?�48�8�Ϟ"�F��Jڟ�I�9�;�0��<�湀���q!)�#?*��{�?���t�/��
���ZӜ`p7�ݝko���^]y�
W�����Ix��Eф����;��;鵉~����������+���;�d�Vx�@�/��lɽ�l�����<w����ߠ�w�sh������A b=�}y���J1RtvsY'p+�F`b��� |sh ��T�0ӄ�@��8�b�:��wtuz�
�ר>��K(��^���aPT�� �D�-�Ko��Uy�*
b釆���������81 ��3�-�!x2`!u�#�|� !Pm�yĬ<*�Ά H'#B H:#Q�	(�UwB��p�(.Gh(Hj%�����E�sV����ABѶ���h��i
b����~��g���*�����\����"oJ����A�g!��$6���������E�w��18f�\ľ�����S�c�����& N�##̆�����_�+9�+���{bthi񏻱3P�^��f�W@�%��i�����e�Ub_��ս�=�B�KG�=�/Ɂ�S?������7�2��'��w��Y��uQA_���Q�Q�3#iݻ-`�� �gwR����ր�_��	�ڴz'`p�R��u�w�c�n�b�cw�[����hbF�����)�ֈ�t����A�+ڗ9x,c�}�F�-��C���һ�a�u�*�)j�����'�҇✔����N�S�Q� ��o	�E8gb�O����^�M���ڈ��me��'wS�r��T�=�G��U�V^s?�&���Ĳ^]��TwQ6;�lkxrxʷ$���,ψ�d�g����s������x��p���dz&�,6u�Ʒ�_.܍�?�ks����HP�����f5{t�"/��Iѣ�*�XL��R%��ݵX�Fh����n	�%��O�r2��9�5I(���LΣTQ���	�*���Y�t��*h��:��B,Z�;�����?���M�����ó�V8��k��8}c�W���a��=����|�����zy��b����@����k�5�:H�T�P�{��:ߣ�]\�?�q�*���`��0����C���һ�1�_��J�.G��,W,�Z���! U�/��n�Q?���P��&Z���F�<']�qZ�⻩lrs;�]��K{:���0��;���0�j�ꯇ787(dXg��@�a=���'�A�����#rHLtF/i��Eے���W�C���=I�eKhd1�'b��laRֲp2U�����������t��g�����U������L��j!0��-��F�QA>����X�<kBm�U�C=2Xu�{"�(!��ԙ��j@
�l����
�{�	� ���B��/��E�����"��%���V}��o~8���j�`vi~9ʧ�%K�@)n�ל�V���X������|�2����z�-����Q�x�Qrc��^ި���JP�iR�E�4����D��C���\D��r.�JTK�/8i[�#��xSQ4 h�S�	d�`�?7'�N�SB� $ w�����_<�
+5���c+ٖ�5�z'eT=I��f5�KN��M\��ʢ�H��@�x��p�dr˪��~��P	@���v�6��3"�p���h�v��$�L�x7V>-�q�ѕ'`k�؁����`<�S�- cE;=�T�w�[N�kC��:~��(��Бc}Ađ4f6\\�4�u"<Sޕ����<�]�~&��[���U����GM��4��v8�w��ȼ:6v_�Ӄ8b�[Gy�WUI ���]/W[z���fBծ�`R1{����ǅ��G�o4Uo�-���Ԇ^�ʭ��1v" o������$�`��/j���y(���hC�Oƞ���߻�#�
ؤ΁S��e�g�^�u�C9
e�0V���XH����up�Y���!��4<F��}����+��op��_6�3' �N��c�<�=1�4�8������Ҭn�6���Q!�d��C�Ű��d�ISBMNl�Ti�|l(�̊q^��:�����a�T�y�=��Z���:%�%\�V�<����@6`%�~�(MG|�J�L�γ�Xs��!3[-�O�U�v�,�<�[�cv��e(�"�F�^����/+@y�]T�-WL�5�׆�mm��׃��N�M��PvDSl��8:'�Y�&�v�n��Y�e�'��M��s莰j���n���p����0�����$�u��h�����k�ڄu��i���\"�������Շ)^��X�4.�U)J��W��$8�ڝ��V�,�
e��~����6�f^w|�$1V#�	u�J8�.��R�Uu�a;�a��"]ƈ��#�,�~-.�Kkhi�*�w3[U�l���"�!��g��0Eo(U���Aw�����H}v���<&�:�����H���J<|Rb*�ӄ6l(���!l�M�X��=z�|�����m��ч��4e�:ǳ��8��~X��]�� ��&y���1	#��?��dr�����!��s*��Wv�d��G�B���İ�^�NDow�m7S�R����Bm�I*�D"Ԙ8�OrN `�d�Yڂ�4��#J��eGq�q�wT�p�x"�3���;�n%�����庶�V�,�*Z�dZ�o*͎I�k���oB,ܝ���텱X��ص���� �,u�r�Л �����i�55@8
"����k>\�S?��S�����!�N�3?v��@㿫��Tȯ�8�,.Z��S1�;��wA�Tj%Vgf�uP�BR��r��<[�%:F8qG��#�3���
֕��ED2^�ib�� �Y#�I�A��ш�u@M-9�6�~¬GG�bō
��7��zԁĪS'ʪ1�%�e����N�+M��4o�o�{����ƨ5�ɉ��/��fa*���F�c[GVT�����ϱ���F�]�bZ�$�Jͺ�>�n՗��Jz}��Z�DD���[:S�� q�ԕ�*/��O��"YJ��#�z������R4X������^Ȳ�i|���<��6nJɉ䜠�i�a�eh.���XN��&���Ud�1��h��䷷�yG�P�W����\�'�Fc���ͅ������;�3�ȋ��$}�0f�쀚Uik�s��8�v����q��6�WA��Xy�HŚ��+��=��HK���{�uĥ����aI�Wѷ>�V%S����Q����Rπ��1�}��b1��t�E�7X�_u+��p�xF���p�7�C=��sA��8,�~r�-��.�ᵣ�Q�Q�s����gp��w��&���vld�0��oN�!D�N����g�T�����6��#��>J�ɔ�%� f?��dT��\s�oI�_��c��>9�F4��;��ҝ#�H�B�,{��)��R�3�e�s�צ<N���ˋ`�=�]K��}�Q7lx-����6��/$���~� Z$6�#����
�LU��"�o؄�g�|�LL$A�\+��H��
vw����H)�#"���N�T�?טkܔ�(�m�=��1���"��
x��No+�됮r���(��~Y{����$��/2��@�a@�C�rj����x���L���Ѵ����.�5�,�5$�=��c��|�ZK�I��m���e�M=����_��j;K_��(A����cR�����{~x3��S*J�{~�;#�S������˅�	�]\�kyB71ܫ����Wf��nz@�q�_�mdq��ILǦ��M]���a0����$;=#��yǶG����m��b�����6�Tk����ud�o�_�G�| ���UB�
�uQiB./'�SX�H��gRd P�Q��! �`1�����q��
�}.����:ٮ�A�������^=��&��&�V�瞡º�RE43�����Ž�ڥ"����za�"�����M�Rd�s؃�i��6�s�"���k��E%�1�	��I�``�}C](Ki���vR�γ8�柉b�ƨ`�]�F�a��ȑ7E�8c#�b��)��C��`W�K616�X���K���~9�&g=>}��N{Nz=�� ��%'�0�+�A"d��|3Q�]I,�j�6�u�`�f��J\�)d�fѨ�a�!��{cz�;�#`Q}�,u.���g���F�w�v$׎Ÿ��W�U�2��K}y&�$,V���C��]��4r����$�!z�Ʃ�7b�8'[���3�i[Z�6ذ�Utn�YK��*�LTIB�G{8��@Q���>R�eR�^� � G`AR�{YQ�M2͙���$O�'���L��3����gê���Q�����_ܚJ���z�M��)אJ���~��,�v�!
>����T�Tl鱵���)���&�z�Jvn���3(ik���~/&ւc�����#�xt@W�s��)�����#�q
�W�S��+=ϰ�&q��^ 2�N��5{�4K(�>���p%͉�y��aHJh�2�A@��Jy�Z x�+�c�'�vz'���t���忬��n>&�� ���љbz����2�3(��3^w�|b��*�eO!NC�T��i�b��2�}�c�{SЅE�
Ɏ�gn!&�P^�uc�����&"K��đ��z��p!���@Z������M݈M��+R�L���A��pk���a
:�3H�'h��4yl$��\	]���s�	�|q����](���j:T���nL;;�며����gJ�GN�cyS��a3���Q�^b<��9p�}Y`����U�`���?�WL�?9�h�P�e
X�\�&GVg�^��1*5<;�lh�5�D&�l3�����E�k���,�6�l����7���fU\^�����c���톇Boig��,�vX�M����QB���q�3,j��g�qd��G���鈧XN��k�o�֦�mz�d�����z:�~H�Ʈ U�o�&��QiQ;_8R-���޻I���tc#j\'��GV�wΠ�+�CӁ𰙞�g�H4O�8��P�&�Hk�gX��	wv��Y�{Q���ӳ~��F_M3�� q����OVI��"á;�|'��m��V���"�`������Ɛ�����=�i���ŐZ Mvݿ-���Ŷ�
�.�Ȫ�����lsO�Ls?�E֥^ۧ7����#����!�������Lw��q��O�M�7FP�C����=6��v�i�r�+��KmĖ�zP�'��d�wU�D�)8�<��H�Jr�/�`��6�{w*
o���ͥz��|2��f��:X��k;�ʶa�EV}��B�?t��MY��A�wf����Zr�����)�*6U8��t+�L5e�_�)e�ꐆ���K�\W-q�)qR�����W��v6(����u�w�v-�����Z��L	sZ�5��@s�>�9޴�s����f,�@c:�������ٗ:g��}BK�=W��
B����C���wU�l�z�1��� ��%��Go�����hB��1s*&�4܋u�f�)7�*��N��䷑Y@��{Ι*�#fi��x!��ʊivj�Oψ@a%<\�>Ɠ-V0�[�x�A/^0��4���Ka`N��Q�3(�=�ڐ{�z1�S%9S�ly#$�"��f1u�V��&n�Y������7�#IߏV�8�[�ԏN�S�5U��)�`�ڛ+���q��ݿY�P~Mw�J&����Bo�d��<�d@����8Bc�B�@ba��|���2��'��F��M�@�܋�E�Q\�Hư�("