c�����V��������`�7�O����$��"۾�l�k��z5��?�|�
�!
LP�m�&x7��3�����=4F�@�`�n;�p�mF���ĥ�Vz�X�5^H�%L��@���MjK�=��7�Q���Q����.�Z�a��ode�`��E����P�:�n'I�¾5���i$1Z7�gwchm1��B�N�L��y DM������Dc�܏�v����-�$���Y@k�g��W+�\��#�F�b6��L��'C�o�J8�ք����g����D��C�����W�'���̛�@�|&���
��L�ʿyī���>m(���ʹM'�� dޠ	`>'k�1MQ�Cx5���^�p�<��1j7�.���r`�r[ޔ"Lw���Xr"s�� o�T�\g�kA�u���0���za��SM���+ʚX���k#،h�=�&y�QL��$F�qH,tQ�3��,�A���B�h���^Pā�5�t=��\Ξ:!�+�p.�%@݃���}4Q�ۓ.[:⩑sx�Be�H��b��О���Yz����S��/74'��"=�
)VY�>l7�#��<�Y�:�0-�b}��x�u�������x��~C|��u�NN�.��!�2��`�M�r��G3���a��H��nB�;0��Ԝlo{��|g��<�fBÀ�ݒ��q�>�jdL@Ԭ�~��⢺+S!�ezI���\I�o�����zY��PB���˽��I4C�LB�u�v�mn&�Gw�]^�*8D�O|Q��e�.j-TvO4�Q�U�v�|�ɺ�Q������{&���qt�y��9&��l��	��şJIi�������t����l�,�mo,�O��:i:�����3^�8�^��u�2�p��?g�ƚ���a�]����i}������!�sT
��k@.����n$��	��f�R�"���-$8��~��C��-}�v��nL�4�Y��)��Lg�X8�T�iX��q����8k��A1�/h�R�������T�����@�[�P�Z��v��5,��X'lb;ҷ��������£b����"
����\���*D��ȣd��0��1�����e�DC�[�����D��f��M��̐ۢ(����'�!���2��b7g?s�7`�e�Y�<�{`����0_`��Ęl�᝗CHzx�J�-�$X,�6 �(m]�[�
�����F6��~o��cX����I�@L1P�zN	>�G3��<H��F��pc��y<�𚛊Y�Q1i&�S�x0Ύ���f1�q��C=�x�0��Y�����s��{�Q���Up� �Ʃe�_�+X���b�7Ԭu�ު�pԺ��@���N�O��~ܕW���9�6���7b��}�$�k=���>�S�_��h<I�ml��;���1_�\�ADQo���ڏ�;3����.m�wVp<=��nc�^5�Cjx�1��4 ���O�Ԡ��ST�ix{||�&}�C��`�9���=�րL�w��Ū�ő����\-��50>v[�+hq��	��P��v�p%������h��x؎=v�}��?�M	���RdT4S]��Uޕz{pDE�<�7�����oL�N�rJzJszK e�T~Mv�-���ǈ�\���i��g~�-x���}9���Ý� _a��q�^�9�3����iW�	Pr�=�Q�Ki�}h@��\ܟ�2a��!�	�ٿ����;���V��� �����aYsX	���sH�'�?��Q���#��j0�	���e�x9���b��顚������."�����r8h����~ґ�����]�'�Yb�^���%�X��zAU��^]c�3��_��