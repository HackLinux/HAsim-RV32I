��g��LDK����ӧ��t� g��ic��2����,W����r�F�&#s��L�B�S��,�dL7���d�Vs7SL�Y?Tꇨx�Ul�;�:�AgK���B{Rj���
�TS��:�e�T���
����i�5~F������|�&��N�Y���eu���ea9ž���	{�W��T�:�\<�f�|��8t�[bj�E�ɖ�rwMtj&�q���Q��5�>�ʵ���s��y�\�1�a.������,'�cGt��zNI�爅���b���e��)W���8	�g&U �]j���X��*����sB�,�|���U��K���_7�j�R��w�j���H�p[:��_���v�	���a�Ø�Y��8ٳ�k�S�K�cgy�z"b�Z=F��`�QS$K���Z
E
D��w�?˜����֙k"S��P\ F�Rqzw���D�~��#{��L�F�T�F1��k�W�`LV��u�R�y*�)��hzj��kt=*#n�(�9"�,nr�cՍ\�^K�,��u\��p��#��z���g˒���3�O�,.>��fq�=P�֊n}���ޓ�<wb��>��0�{���DkU��?I���Sto��9mǙ�yS��lǚ�yX
]=;�S���-V��!}m}漟 ����ko�O�^�����u�O4u�v�%~�ɦ&�ܡ��"g~�:cZ���S�ދk�s��6d9T�wǄ�lD�_E�������eN�.�V�	��@��J�W�~
V�d��B��V��N܆��P��!Z7D��"�^&�	Ӆ��Q����}&uv	a/2�{���ak3T�Cس���"]����[�k%��Ӑ���r"ow���_��g��P7����Q�)�x���g�?�=�L��������R�[��g��J�����r���=��I����bt� ����I�}��Z�{�C��B�z�L�h����W�NdUZ�Up��2Q�L�{�E����{��?iAG�����J�
���B���N7�K��8��N�n{S�*,��W����8�U~H�����e�܌���u�U�	�{H/n�{���z)��j�'��l��ڇ,���%�駍�S���z� |�?{����D�nB�Uu�}�UC[C�ce���:���g�U�:{O��W��������&��y<E���Rt�(E��RT��LP���R���pm�i�!�{e����JV��g{�v�|+��*�ޛk0&ԙq���?z���p�Tر�����l��q-��J)��(�K���^"�"a��^"�冎�T����tj�'R��h�{z�V��*�q/Qu4u�^��%��!.t�FZ �z�V=EEEO�԰����XqU�HL� nt�o/��5�:=�r=$��������@��Pړ��<�p�)�]������-}&i���>3��:k�Gz1����XO;���A�Ƀ{����О��T�Ҷ�̶���Y�o��R������r�!&���Q���*-旧7����^���ڤ��CTA�����7�����-V�K������Cc����C����7N���j�v�1�~0�ֿ���S�����^�����{�w��u��/�=��B��r� N��=��c0��I_ݕ4�+��#�Q��{��Y��l�O�3ob~�^�S��G���+��z��ͼ�E�J�6��p������̷�n��ꌶ����I��xS�7V�:K��S7z�ܞ��|�X�JZ'Q��ڂ���@�y�GPPu*�˩�3�S�U�Q?��J�;��~R�����W��=����B�Z)k��p}�9��(����F�gI�������R��q�L)ǩ��KI��͞+�+p:�Ө�%�A ��� �}2��]F�:��é�s*aNA�G9ϡ�ۢ=p!���bl�U���,'q���aj����"����g����yF�kl}VQ��Ĺ��7R'��7aC���\k���`�?lU������;l}�P7}��~^�����vL�>����!�YGR��X_pw@~���P�l�+T��ĥ��p[��R����R�ou�_�꜍v�H�Z[�z�Zںv퍾���d};D�ћ=��<�uFG��ZM�R�Kȣ�C�W��g[�3���i��R���<��X�[�������,�x��E�EVB�rC�a� Ё)HG��T�a�u]�zғ>�o�a�D�s�ھ�_}E��d�\J?x��OY	/����W�g�N��E�חH�d������ڡ[�u[�W�]���m{��`k�+�oS.��wis�K�!���������U|I[}`��ڔ��Om}6PR��S�5����|�5��aC������?s�	��k��~#?��JB���t���ކTg�t�b�Q�=X�,ڶ'�z[o��W!�y9�ͱ��r�'��>=��7��*�ܺ�>o��o�PUn���l�c���L�穂J�"l'�9�a�A�y�v榎�O.aޭ�Q�wm�>�:�z��U)��6)^e����E���gU���gԙ��a���0�v"SP���:P�e��(�n`OqmX�S<��8�k��G�Vqu.
�F�V5��c��]��qM�A�c��!�Z h��Z�h��=�y*]�RֈZ���jm`�^��P�|);�	���NVL=>�[Tv�U�5�"�N�y:ź�~��~cס~c�L5�_�J>�|��ti�����л�-C]d��R�����%�?b����� ?�D��>ûs_�c�kt�P�F���CKO��y����ԩ���d�n�Zzk���ﱇH�"[2|�Z�1k�!��ꥆyq$᪉SE���Q�n��o����1��b}��2�ª�Ice/�?�m�2'A�	̝̟UX�<9�v��:7�>6��~�jkS�á~3�J��n��bʸne���N�R�)�M�]A\hc�U�L���� ����\��/i�f�v��6��U��m��]̝�̝�l���s�s�w��Ӂ9��m`�z�3��e��.��i����G��Q'�9չ�j߉�bϩεH�T�'t�TgT��Tg�^ȘP�8d;�.�-Nb�G�A��6��l��e��I�+T.G����"�����N�ﴞ�7��g�Կ��l�sW5�q8�пC�¯�,�S�MRy �u�I�p�
���m;�pP�c���������T�=%�]���i�}�����7�7ަlo�_�E����1�����\���i�7)�����~I��*�Hh���\����B߂U���v1sz�8����ҿ�踙�	]���ǰ^��ޢ� ڎy��k���׷���Y�����]?X��vU��I���v�S����øv5r>���k���v��=�(��(��B�ļ����#t5�g�>�V��9�� ��؋�u�V�*�ZM�![Մ��F�z�X��l%L�juNA}nQ+���V���y�g���%�)��߸����gދI��&��9T�A��7��6��V���j��$y��<��|���kv!������VR��_�����{���ڿ3�2�����p���Ž��o3�;����N����m����[T��?��	u��:�(��I2bn>�873V�W��^��b�ޮzWV��Z��Z+��^ջ��s�]L�S�y��2q�S�캕�����ί����q� /�{����3TF_�^���˝���1{7�(�{�.�7��#]Pﴶq?TνP`a�]�i�=M%�2�3I�{�PyP�t��2�=�:u��Z�g����O�.ꩋ9���D�"Ns��Gw��M�٣
��n�]A|d'tcoG� �l�+U�ån��#�zS�xji�po��G#��zX�`-�E���{���M�u��dR��2�uc��/��>0D���������8��>�/ �{�����ܩWu�Y�ʿҹ�T�D�s�q�y����)���c����$�t�*�{H���.�?�Ŀ�y�]��޽U�ɪ��W�v�.�}N���f�Z�YG��o���;'����M�e���G�g[����ڬ�IP��a�I�q;_�.Y_S/�{
泣H��I��³6��Vu��X���GX����zgV�ת�U�z��A���a9m�W=W$��
�{x��r֗*�f=�`m�d�����*փ sZ
:�e�ª,���p���9���̙�:�^w�M�١����[�h}�5YE��Ӟ�Y_�[E�����\��g��`��J�e�n�����X���\{%����9�.�X&n�W��nR�8f�"��+l=�L� 4�Ip)������R&&�Qp��B�eS	#`.4�qp&<���h���*x��ͧ��p���G`O/�@�:l6�}/���t�	^�/�lf��&�|H�ٰn���>����E`;���M������a��]&��Ca��"8.�����6��C%
�a4B�A\����>� �疉}a0c���
a-|�p���~�`&��Q�·��x��5�>�o��敉>���!P8�!'�9�
n���)x�����#Hv��a8����fX'�yp%����:t���Jk~����0�BX'¹���;�x�������B�eb���0&�L�����p2\��C�|�t�$���!p(�� ̅:Xi8��p1\��3���g�=�v��[Î�'�C�
&�48����"X���t�[�|�A��2�l�� 8�a"̂,��B\�����Z���_�G�L�C�à&�4�!h�$g�Ep�
����Qx��Z� >��`=��2���~�T�0Ӡ� ��Yp\	������ ô7l�` ��aL�y�,��p����x^���S�q��~߷=޶�[��ZysnY:�8F�`��u�+�!-���x�	#�j�d&Zg������1�+�~CCxV~�?x���|�o�P�^q>Z�cL�,�}#����xo�[T��M$<�SF.��Z�@���|E}H��W��]+�'�#,fs����Ck�[]X�EZ�}X{���K�hz�;j��{��ă����(�B*E��|p��U\�%y4SRw]�D>ʸ��n����;d�����Y¦�Cr�g��R�K��1��>����W�ݥ�Ŏ�G̠7���ݛ�[士-���ܶ/B��)V);���؅f�vE���̝�����Y���Xt�T��6�^S\�h��e�����]��Nm�|��ؐ��:ה���5��Ȁ��Jٓ;��l���_����
�F,�{Oi?��[0�^T�,$K@�Q��b�1�`ˣҼ[ܣ[B�3X��;d�۫�E��5������O�N�,9ɇ��
�
VhH�`�_�����Ng��� U��8�_�H����B�8��8�#��0��T� -��&cmխ��v�P��{Q�Vx�s��O�k��������ei;�5K;�$=|���2MH����H�3�HvБ	�]��ti�ĳ�!!��[�C-��� oH>� �?�!Z˴s�: �n�+1^e����
�A�7Sc+e����G2/�l�w+Ɛ����U��sn�Ej�E�d�в�g��DL��=u�r�|�O1��:�������ө����ǰ!hse�ž�E%V]�`�"�$A/�`�צČ4�7 ݊��bf��M�r�7����ͩ?�ck�Fq	����seL�jQ/\'ba�8T������3���~!���T�d=oo��1��$���i����9I��fR��'G���J�<f0}7�1�V'�C�kś������|��[�)��V�iw1�2��&�tf���o�K�C�N�����?9 j������ҋ^�E�+��'9�:�ƅ_�}a29U֍{[A��~L�.U= ɏ`~��^q���������)�X�"�=L�W�R*�TI�@���N	Ŷ��c��e}oz"1Τ���t6�C�����i���mL��f�z���nD" �϶��$NRc�e�@��Ѥ�<�XB�zQ_�4� �`m<�I��&[QL;/�I| �,�{��g��ā�Me5ұ\Ti�NՁ\޳<�'�I�\@�j�c���9�����_�ˣ��ʱ�􈠹��܎)��r�[=�>ԯ�G�9c��9hj�N��"��EN[�E��T}��\���i��AN�\<&�6C�رa�a��a:Ǵ��8�n@\Ǽ�z$���[#�P�~��Tx���������1�z�"���6�)�R�N�+����$��78�����k�ix��aiքi������穳�r�n����</«�6|_�/ O���V�=��0��(�� ��-p4���Yp!��k�&h�{�x^�Wa-��ϡփ<����C�v��aá
�B �@-4@Z�XXg��p�w���8<��{�	|?��`�N��>�=�0��0f�<BB���X��5p+����ކO�[�����~�/���
�aD!98�Ùp>\��mp<
��x>�o���g�/�-a����p���0�P���!�0�%l�C��Do�� �w����([�>bK���Zl#�}�v�b{���Q�$vb�O�*v��=Ğb/�_��}�~bQ)�A� 1X(���b�8H��q�8LT�j1RԈQb�#Ɗqb�� &�Ib��"����&��b��%f�9b�8\�G��b�8RE��:��A4��X(�D\4��H��8J�EFdEN���X$�%�hq�8V'����T�(����rq�8E�*N��3ę�,q�h�s�yb�8_\ .���%�Rq�X).W�U�Jq�X-�׈k�u�zq��Q�$n��[�m�]�.��w�����q��O�/������!������I�xZ<#�ω���E��k���e�xU�&^o�7�[b�x[�#���E��@��������L|.�_�������߉�����G��Y�"֋_�o�w����7i��e�F�����mlf�3�nln��(7�0�[[[��}���;;;;�.F?cWc7cwccOc/��1����������ߨ4����Ɓ�c�1�8�nl�0153��jc�Qc�2Fc���8c�1��hL2&S��F��fL7f3�Y�lc�1�8ܘga�7GA��uF؈Q��h0����h2�F��0�F�8�H#k�#o,2K���c�c���V�c�q���8�Xn�l�b�j�f�n�a�i�e�m����+��������K�K�ˌ�����*�J�*c�q�q�q�q�q�q�q�q�q�q�q�q��n�n�a�˸Ӹ˸۸Ǹ׸ϸ�x�x�x�x�x��053�m<n<a<i<e<m<c<k<g<o�`�h�dtk���W�W�׌׍7�7�������;ƻ�{��F������������������������������6�3�7�c�`����������Xo�j�f�n�a���7�����-{Ȟ���-7�e�o��rs�Y.��}�r+���Fn+����?��r���I�,+�.���U�&w�{�=�^�� ����}�~rY)�A� 9X(�ȡr�<H���y�<LV�j9R��Qr�#��qr�� '�Ir��"�ʀ�&��r��%g�9r�<\ΓG��r�<Re��:����A6ʘ\(�d\6˄Lʔ<J�eFfeN�ȼ\$�%�hy�<V'�����T�(�ɓ�ry�<E�*O���3��,y�l���s�yr�<_^ /�ɋ�%�Ry�\)/�W�U�Jy�\-���	t�q  p��z�ܷr�+1���眳�ܥ!���y��ØU������Ծ�����!��c�<�ߣf��o����jӢ��+�C�9�RA�NÆ���M���[k����I��Fyf�#��;�u%��H��ڮ�E���3�]�,�\�.:/v)rYVS�{xp�}l肼�\Ï�.��
e�W��]Ϟu�U�Uˎ��i��?<���Ʋ�ZnT�S��h*e��͊�c�?��W��C5�QF���x�b��1�����P$WL4:��b�
�=yr��:�.P�J0"�%���oe/�|\c�Z5V�:W�Uk�R�Q�Dvt�ݙ���6榎��2s�P��l�oRK?�~?=��=Y7�꣸<��o�y�k�'�-���4�{m�rN4Ia��&qM��'�#���(�O�M�^K�J�D���Ym�(û��y\�ݛ���i&�F+E>g.o�ؔ�������-̝̭LS̔����%TWj;Z���m�^�'�}�=^�G�T#5��t�����oȅ��;�ۄ��-B�P����-�N�N�N�O�S2��
;�T_g_J��Q���;�X�;��:ڀ��dC��_�e�9ȁ�2c�c�19ރ��Ex��ޘ���t���C���[��-v�]d�e�l�ط�9�ɡ�!Nhb�ku2�i(-@��Cb��DW�:�A\d�c�c����(%�J��Tx������zv\ʑ�rv6��6��dM7\�����g�w�+$I�#�*����i#3�[d6i\��nK�QI*�J3]Hц߂�F����/�Xv�S���Oj���;@���6�N��q��M��8\V�)�#;g,t�����J+m	$p��ǭ�N�P��p�3<(;�v�{����V|�8ٝ�J��{�׎6jG�v�����<2$����p���2їX�]�A)��0���W�lP��� J��j z�ui���i7��!�3�K�����ɗlصa3a��ɂuO����y�.���
�)f��W�`X�V`%�@M�A�hZ� �X :�W�ǇC��
��j��* ����$�Y��^��T��Z�P�U|�m�m�Mf��i<VJ0�,�E$�$�T	 �( �ȉ]�iauxd�#��y�F� ��C�K���������$��_��N�"�~�����nLd&�C'Ӑ�L�����y4Mw����i���Lue�*H����;X�M�(l45>j$���QuG��f��C7g�dJF�!���?82'2��i�1%��"o�^j0�Ŕ'�}ّ2���a��{^w]oz�:g����J�a��]�׵�/*���9���M����澑��D	E����Tv��uC���,q��Z_��g"��.��^����k���Biގc�᪟��![��kf�UM�����ZL�wjGt�&�Z:���}���֐��?��pmU�۪��U����R�r��l���t����Czuܾ�R�Q�6�������a76\;]2�i���O��kc�s�A/��Ɵ��%������M��|�E�*�(-��r��6���GE��I�uP��Ձ��s��J���B�q��j�����4�*��o܄jÖ�T�MT�&��ƪNѾ��A��38�/�7dd��.-���Ͼg/fw&�1W�\�@�φU���*m=���|������!�B�h��j�Ux�=��Q=+,xR�hUUiܠ>m ��$2�`�d���T6g�T����?����ы��\��^=.0�:8a���g�s�ȹ�K���	�_��s�p(�ИZ��D8���2�h"�XE�-��E�L��T�r�~�����N+c�bJ��������ʦkp�ܚс��N	���2s��n%&TKxU�R��H��i��l�d*��a�8�W�G����|�9�E�:��>�4D�N��ڞ�f�*�����deռ�`�ԋ��v�t(���T�q���?���"��/�i��r��n�n�1���S
�qS�g64k{]�>��nت��8=^u�����KepӍDޝ�*7H�;��`���+��KD��W��M�ޔg1zIںFK�kS�1���h,�1X3}fp�̚��)�g����tBP�W(�Y�hfc:�/�T@U'"��X�I������PCt$��v�H��HhqF+��D��Q��5P��;Z�g
�qԘ�u�~�FDpF�Ufl|��t}V���Ne�#������\&����⑚P6��۱�i\4��ak�*8V{�BS��PK5��{�Ψh|#b#�&l3�zv4\4����?�3�(�c��(mԍ1���Rˠ�M8&}ZH!E}���O�6�)>�A�8�����m�g7��Ww�X���Ic��b����A�����	�w�/�����E�s�b:M,����lPg̜>~�ؙS'�*q'�T��du�`<3'��7�zַ�-��S~���Ks]0�K�C�6e���f"���XK1r.ѐ�#�HP��V�E"^�P��-6?�dL��`8%�Ӛ:�yWЃ7wNgR��ml���68xʳ��Ҷ�c�6��a����`c2ل�����Pj<�dʊi=����	U�H&[1��u�a�>��qf|N��:�-����P*�+�u��s�JÐ/��ufK��!��t��E,�>(� ���Z&�	e±�����^k��-�U��ǚ���ˉ:��u3�'����9�.�#,tWmq�b�S�MD����K�͑x�՛��M���N67;U�*iɔ��pD���G}1
�(�u��͡T���d&Ee���<w��PS�`���Tֳ�}j�_B�r]KzQRz�W�|I�����d��%|�B�ū�+z�!U�nV
�X��T夣�$��!S��si��Li�8]��������1X�C�F��2dӉpB�C&�b�e�j�,fs�N�czjT��>��,�1ǩ'M_�e�^/�`.1jJ�6zQQ/��1���R�=��1@���ʢ�8�T���X쬡�̐���>�˕A�9R���J��&Ȕ�+���>;������s&��Usl�5S����7��(�/Hs�!�L���W2����=t�zOƳ�t-1]ZzWzq�^rq7�:u\���s*�ߡ�����h&JsX��&��;ӘT����*�3g���hɰZ�� 4h�AW���4Fbi-Һ�2�\A�W�N�9R�eiLק��-Փ���7y1�����z+66��aC�N�Su���b7��r��肢j�SS>�o��TǞ�Ձе�Vn��΄C��Z�h��)jڪ���
��W�jDWѶ|HWJ�P ��,�)�^��뎏��|1��b�L���^Ã)o;���{%�t�s��z�*�4�\Jҟ��:�pK��ԮDi�;L��q�xݿ���_X�I���K����+��Ly�5���s�<����Cc��z�9�Ug�yΐ�T�.@�[����F֫�.��)au����������굌ƣ	:�_׳�r��ճ�qG�R�Չ��|7�������˖�x�Y�{���=���8�Vvj����p<��yWQaR�([?='֧ԉ������b7����zǭgܹ5�F��.���Q]���s�F��?�#�
ϓ2��E�o(�bD��)+�Se���r{B&r��Q���>ũ�l4/�W.'�����W_�3
#��8g�3j�1S�(W��+�M ��	��d�/�4���!c1#ũ��?_4�1���	��/�K7��W���]�������ݞ���(k��GR��g(�d��ڿ�u�-����٠s6�c�v�Zw�'�'vú9g�Pz�L]����
�#���d�u6u����J09��.�s9�`�U(Aޗ_u�E��+��s޹Pį�Db�&g��t�4������Ͻw��e���)��bN���#��:O����|��Ηf<��<�A��W����~O+Z�H�4eU��"8J���Q�XG�3�R�һ����`��T2�
f:�+;rO�������0��+Eu�����;�&Lٹ��'�e��ͨ�P߸q�O�ՀTj�1���b%٭��ɽs��5Ĳ�ڐ���ZD�%]W2O&��\W�/��}>\ݯ|t�~����O��4��P"�