`����W��}��Y{��ݟ�}�s�����' ��'F�\�9|�r����,���~
�4.s�q꘸�7�[�7�6c��E4�i���Ȩb1Cr\|"���A۷Y�>�b"��|xJ���>����]x2�w�ԥ��NZ�a���C�E�˪��[}�
���A9y;;�O���3�c;u^��nY������'(ty:<^�
��:�z`��2���5�:9O� %-Y�J��
�F�%ui��J�Fe�&����QG��{�{,�v��J�ю|_�TXy~�e_�ѼKnkjX�.��[v+#���KJ%N����8�����u����|���H.�ӘlZhy3�6��8�������	��n'�_�L9��=ƨB�8sX�Wf�r���9eIɝZk�t{̢��5��s}���y�[�\%����& ^/jl�>_I>�������QhųŖ�Ie_���~�U�T�F/.�������MQ+�Uy�}��^`���?��tGRa��8:�`a����3�9�watŪ�k���'4���"�@���֚~�y\N��י�i�2kg�+�F�([�=E&��5Ä��*����ʷG)�\"��=R�������?�y�
�]I��;\Nr��E6�~(����&�#�;��Ztt��S>����
ƭ��y�����|Xr������N��̻��W�a[�^B�:'~	�����0s�ʓ6E�]p����v!���&�Nhb���!�%��tF�T��\�nTD�a���Ce[��_�\��g�	��G%4��� }�]����������dX�lɄ�d$���L����$3�����G�%h�8H���<�-�e���R4Jޕ.��0;��z��a9*�;�c:�:I�A��{�&ODB_gL�'J���-��l\]v���1�@H�6V�8sъNQZ��|���&���b#A��M��bϕ�w�C�чп��P�9��vG�H˛<߂�Ns��|�$���3a��'A�o�F����;��`��@@\0�'x
_X�4�Dhq��ׁ����߱�>#��ч�<���EܭPl8�g�9����5��Bi7ش䤱ݛ��5�䜜=�l�Q\l:�tYX%:�G1�b���q`1eճMA&F�y�s��Y�7��ܕ���g$Z,��67�"^�<��K��1���1Os$ocy�b�tw��P��kũ�d�3�滦h��>�Ҿ���ۍ���n9a���m��ǼMx�����
?�;��a.;�'W�2�JVb�GbP&	�˛N�/���']Q2Bw�;������d$q$��D�~��W|5,���)���+ӌ����PE�K�6eӧޒwv)Bm,هEgd��_�/��{u�����?? �.	�`��'��Ev���{_5�O��%������e3c7ԏ1!X��ϋ���M��ړ�W�}�*�JN��\sBC��,N���>QH���$g*5���d��^sf��e���y[e��?is%�wm�G~Xwqy ��>J��.�ݴ�H
~�[uY,�U���M��'U-6�����}����-������� n�]J�R���t�tī��_�v*c>8
 ӈ�@d���/��-o?Fo+��*������^$D[�G��~[F4M��N�[�D��)��*X$���1�e��U���E��3O���@SU1v��yˎ zN���bk���X>�p���� ����mhȕ�"���!�Y��`��w�;��z�S̗jd��%Fh��i���.]����ꣳ��?ɥ��^|쐺d��k)���4,�Px�]���O��G|@��8<{�f`��zM���̊k�)��B��fcK�|:Κ(� ^WQ��W31y�Oz���W�C=��d�wř�i
�� [#�nZ0c�;Ui�H!�Wc�|!�@�H��mc�����*�xd�jՋ̧Ϯq���pG���w���5C�J�H̹�42;��v���Bo8�b��;n��}EJ��|���E�4.�*x�]��$��� u�~��:�-|�^�RǗ�W][��T�^/E���A\DA��ԽX�d�zc#��Ӂ��i��
�z�o���˿��@�?���}�!��x��~N%C��CNRgϱ���x���
��s�R���������8Ø���"�V`�@�� �c�)b�����������~F�R��/�*��Ӊ�\��of��tQ���Uc|7��dx.}V-Ë��e��avdդ#��#]�����E���?��?�Z�:��UL���K�5����~G�P|aI���׷�'I1��@Fm��&�x� D�c��d���Z\��Hr�U��yp=J���;�.�UiS��P�AZ��r(�]R|޾.s���T+x@�7'X�I{&��,A((�W4C�~<�|&��eJ<��GfX���e��k�ywɈ���):@r5��,�&��O<��!�=B�L����k*�QS���5�.\�好���gK�O�8㥡���wp���{���4V���"��}���y��&��Q���L�s<�w�#�~�[��k�3A�����r��:�`G&K�