��B�Y�^��X�Օ;D�`	yAe��g���8�
��59/k��#m�)�-}ŬR��,tA�joj<����HP�U�-��G�>9�.��f,<���(�}r?$2^e��	J�ł�(Ч_�XqfPmvh#|���چؽ�O��$7�1��� �E��C��;��I6�����}bGu�M�͢�|�)��C}��߼
[������X9KdH=^��:�F_@�$Y���ҷ��X�n�i��xż�3���$�ij�]�k&4�	�{<�V.)h�b{[ �䮼z!��N�Y@(w�L���j�ntzl�uo�8�iU8����WD�M��,����(�HJ.�����
�|sIV����������8j�aGO�ї�$��|��g�.#2��$��,�xq9�e���<%�0G{E-�� W%���m_N�Y�T�2���^#�
�sq!�E���}�s�HH��|���K�Jv��PF����ړ�LT��sq��d��J@�t�- �����$^���O��,~>�8{\��L��{S%�}����{��j�`8U�����퉰8�3�w�>5�p-~N�)� �zL��oR��I�YӞ�<�X_x�I���2�&��}�f��9��M+�N'�$MƎh3�v j�q8ahn��`^�h晿�O�����PؓQ�*��Ĕ���BG�;�5W��2�y����B`�I�(��M3��)d�6]�,�Z����q]�ԓ]ZJ[�*�"���$b@�T`�E6�)��ݶFΔ])�rJ�d(��v`�*����}�Ί"��A�����̗/9�G�������2XI�:S���JK0�Ek՚�r�\�U����,F��7A%Ų0PZ �]���;Zi����+.� b����T$��d���|�d��M���k� .���2g�k����w=�p��OU�#�IK�B�ϳ(?�-���5-�^�&�u�/O�p�fK�mc z�|���.TP����8����k�d�p�y�"��%��%�Tc��:�4)R��r����Wc._H+Ch� 焽��Ͷ����/Z�R�i-$pjԖ6�IfN"R>�H��������y`yqK]��~�,�\�T����:�>]�a5�}σh�ꀚ�;1L�/�ud����2�	����-��"��V�yksVGɸ�:�{bu�m�D��梘�2A+�64[�4Mi��z|�.����kJ�V��Jdb(�l���j��{�J�:xKix�hKQ}��|�?s�j[��X�6�K��e'Tǥ4�4�ps���K�+8����Y����q�Y�d�E��Ҋ�@@)�E��E�	t���TW�K�Rf�!�暵�R�/��qe_|�r}�+D=�����8��d@�AnT����x�#B5 5�)�ɰ���|�"�1"1��X�O�?`�&����]hZ�"�kK��u���&����M]����j&�p���x�&ؕ���ս��[)��uǵP4�k�����= �&)�O�3S�8hh:ܜQxg� ��c�����	�a�y9i�0"^�����N���I��Z�yڅ{_��FW�	�t"�M�~�k��D���ݬ{E�Gg��@z�*f��]c��n:���]h� �J���uq�!���ұ����P]wʸo�jgG�����v�	�r�t��Uww�8O���3�gU7���-'<���No�gz�6\T\p�C����'Rf���!6��5�&As���d�y3�i*��r���S*����Wka�����ȍ�I��!���������P
*��*�t
�0M�������϶��@��6�{��*��t�DR�O6f�X���'e3B��~Ȯ��m��m;��������v��~�0�
����G�,
�C"]vB�e�r��bL*	��|�U�WM[�<���d*�
Yw���P	�"X;�⊥�G`$"�hC)�~�:��aQ�<!�x�==ԣ0���E]lnu��'L.�Q������?"�~�$l��yq!Z,����^�/@��\�vv&��Z��a�f
�g)3���W_�w����xŀK&t��Ź�צ,Ե��)��CG3�@�>� ���G����H��;�wWy)�����;b�&���E������#����Ge�Ť&"Q>���}{3�	TR=Po_�m{��X�2�����,%�VIr�K�����7�|"hL��G*;(�[����Tt܉����/�1�Z�#W�`/Xę!�s�ϔ���#QV-r��&^<�[��9!q �A.��?T=p�/��s��.��~�a��_4CP�먱O�I&N�1�hU�鏆Fi��~ī��2W&�����iG:�����\h�f�mXʏ�BY�,K��D\�(K��*���qC6��T!��vƵ���TR��g@�Gne��M
OKSZH���`��k�"K��LR<Gwݭoh|F>�>2�P'�)F9�D��u�S	/�%�x�$�yE��1��|(%�4^���XԜ���|�>��O$[-�y{yzX���1O����Tb'�j@�i����<kj`�*w����ҙ�T��6�?�Y��q+XY�,�8����gLiV�����p��h��z���_�R�z�O����nÕ.-���N�����&jO#���[�Y��R������Z:6¡��4+�Ityr�ݖ�Αc�(o�@��#1��ۮ-�ɎU�{5$
����z��)�q�f�����k��W c����x4���Q�r�A��(��,��T�\ 㨼���#�S�[�����s"ޝ�������O�yW/>7�U9�(c��B�܊��'��-Q�u�m�7�B16,yP�M����&"�Vjo�A"7��&D]�"� �l�����oV!:�&�z-;Eh܉����m��&+�`o��⽋�k��uN�	��&ߞ9V��0�*��$�Ru�GJSؙ�������SP�KN�����/�V6��A��l��vLջ�r+k�sNY{�)���UB��7��z�<{Rf햻n2��.	%�5y[�x�l��t��0G���B�&r'`���`���@��D"D�&�������a]5����Ë	�ϼ��y��߭��i��K^��P�z$�n�)�i�-4.�0�����D5�����6+g?���	���,AN�>6��k:L��HHh�qi:�����cuڃ���p���a�~�OP�*�'�B���W���T�B��9Ym������\�MK�E+5gѮ]Ki5[���v�J]� �ZDV�drj2��Xt�:t��\I����D,��)!V�F��BR9�:�c��[�p���	�^7�$	����X��$�@��K���Kt:���x��H歪�Ezb�6'��Nt�����s���%�K+3��g��]r*�.^�g�"e��_�EW�n7%�����gtjI�Zjo�n1�2��
����=b���{r�?�U+�ÃAI�K��΋k�q���e-�[q_��A����iUWs�|S�e8!w��&J��,K�o��\S:�!n��*�E���<�^�%n�n�-睔�Asc�1�1*�ad���[�jۼ7M/�n�u���":
�U�[�ơ`J��B�+!�nf%�ڕ;���;K1���*�g� ��Uc��N��y�L�F[Owe8��7�:]K?D�,G�᫃-���\X�D�e����S�4��������$��a�Bb�kA�k�;lb(�^���	y��n3r�a:i�E���V?�o�>le�W�g@R�׹���Ǻ-�`g���l\���g�n�5`�~r'r_S��,�Iiŏ�)m
{�{=��ဖ9�
:3���rV�@X���C����r`x���GW�&I�<���B�re1�a���IRԖ�|!�4Ԇ�T��Z��
XZ��p,��]��^���ݱ�R
Y:�Gz,�

�������Ay�-�[v+׵^�Y���a���-9 yA9')��Y���+U��4�-��17󅬃E����0��r?y��Ig�T��K�����cê�F����s�����#0 �-CT���~��8��^�����,F�r���Ysݣ�PmBUH��W���l�H|`��b�^�%�!;�i]7#o�.��Nn�_�I ��A�q� ��H)X�)\&�Bm�2�N�����Z�S�zr��o�˹O���j�9���J�END�6 ���:��7��W�R���l��w2t2��6ງpB�׽�a�* ��`��L݂ٺ�ѝ��xf���Ѳ�U�&�ZɈK�/�2��Jc4܆��fMO�N$Jԡ�;�e�9Ha�W�V]�᝟cN�=�!�ЀS�����c�_!�p���9�I<T�-�%����
@�D!)�1u#�d��WK~��+H�u{{6ɣo�B}�5Q ��~|��{	��/|i���*$k��/�X�X��QU�1;Sn
Q]z��(��i��o<�"�|>e.s��M�+zn�B�yX�Ua^���X����) :��P�2֠$*w�����R�|M�H�`�_�K�Js��X�TA���`S������ُ��0�i�i���(^K��=y;VA��FЕ��xe/�H6n[�I�jw/#���&QP\30�Cp���*Pn���":��|�F�/YDw��(L� �����]�	,�C(�Z�����i�qxu蚷^�tZ�O��7'��R�W�5�����bcl��M�f�Qk�=X��ԥh�8��H�7��j`�M���ʒVű� tEEK���H�Z����/���z�R��Ҡn1��'�31�R���ݰ#���WW#�Ҕ�Ǉ#����@��䥁*�8�k'*���糑�7�7rpa`�+$K:wy�+�#9]��).7��a0nW�w$�k;n�Q���=��A9�p�<������91�0�.��^��#,4�����i���XrM�� �8WW r��e�8onєm�fS��E[� ��&�r[��]7|�qFҡ���ئf-�<��-��d��5��*���.;��gC��"&2��H��̈v�ݔ�����|�V���j�KwK�ڹ��'�a,�Պ0���FZ��@x�v`,H��d�	�� �_��2wVw}u��W�seǩ[s���?߿�$eͻ��rC-bmN�ZW:��'��6;�]2W�s2���Q��9mɥ�7[t�x��'Ȕ�p��^w�<���X�u1��/���A>3�Q`Gh�%���E�,�����A�I�(	�����~�Wg&~_�d+�%D�
�伀�\��y�`�x�8P53o��}��j�?�c�s/�&m*���|w)���{(z�b�t�&栧�'5�m9�<Gk�@u�5��maS|��=�]T��0���`�ܳ�t�"a;�T���Z����I�����C�jz�>�eI_@�X�0Z�����:W�}����z�XE_*�P�8ּ	۵9��g��I�P��-1���[�J'�H�C��nwy�ck׋Bߍ�y_

��t��[姩�˶"�P�~���9e��cۻ��NKG��oTx�����O�_��<+n�+n�3P�MT��6=/�J~�����g�~���7�n�팤���b����чu�W��٥�@���Kjt��J͇NdbJ7~%�8��&��W�cϻ�/���อ/d�S;��X[:j*�γ����x�l?wC�����o���CԵ��U5T��4�V�V��o�d"���X8�����u�/T��i�B���t?�.���st���&t9��O�������˔jѬƫ_�y�����!�"O�%�����64cW����[����%�yO�]W�IФ;��p����ۖ�	 �\�[����9����Z.ݓ��H�ԗŎRX�(|Ӕp�m��=�x:Z9����.��yVt�(��/az?��]���,	�	�|1�J�.��?X�Qx;~"!�]GV�r����25ͩt?8q�^��mͼ�4�7���f�U�$~���"	C���0RO;P�xzeěcA���M|4�z���Q\��^�'��e�q����������T�-g��}%y�6f�F��2��ʦ���*�i	��w�ۓ7���o�"+��3�v�{� ���X���s������/���'Zb�YƁ�3�P�Bf�l�VK����M����x#�Ws����
bF���������Y���K0�.a~tak�n0�=�UT͹�:�Ԟ�+:l>�7�^����AWT�q��,����d��m"��p��%�a>{|g�e�IF�w��Yq��NS/m�*��<Dɗvl`;����`�9V��Y٥��s~���
f�,������"{1
Bpa�"u.g�yY.��w����Y�?�gs����L`�85��M7VT�n�5�x�D��3H�>g�	b�v?#پ� �u��M~M%I��$���R�W�B�9�V����O���ȥ����r��uq��\9���mD�#�����.9b#JD�})9`�:�����-Bo�g�Qx^�.B;�N�=����ZؿM�JL�#NY��	<�?��X���r�Z�ݗ0=*0�H�"nW
�,k)��iݸ!x^j��(e<'��R�Ɖp:������G��*X����f9�Z9H`"��վ�	���-��޿e,��|�Sa�׍eFA!��jW���M��Xt^Ʌ�$��z2/��}��l��э���d�9��(�66����e�,V��Y��_�h-:���0ʓ�tm�pW4�ߣ//�ꍩ��MTb1�BK�2����,�i}�d|-I�,$e��~1A�^[]����K.eҰu�o]�`��x��ReRЪ�mx��)���`�k�C�^}�k����nSG	?��dnE�kE
8���N�&�^�V'uu`Ҿ�B��"3���ԕ^ziԷ�J9Z3��]k���rca��A��X6�?$�����-t��y�"�[�k{���e�_����X����g�	�� ���������zMk����A�%�/-��t�ȓ+G�|j]X	��dZ��,4�BcU�
��o��_����'c�c_���1��H��5�)oa-��ty������w�N�ԑgc�$p=�����)⪪L��>Ox�bvO�������?��iL6�h;@ǟ!ߎpX>E^V7 �;X�4� +'!�z��t�
����f-��oxK4�P�e5s�'�wԫR1�/���|*�,-�~�<a;���o���T&.b`��[S��k���:�1SW��]��L��� ��2ϵ�u���'`�H2��^Fp�ζ3��*����:E �)E�hf�������S��*��(i?r~	��k`i�Y�:�����`��\��^�]��LU�dG��? 	�I}_���$�/'����ő����z(�`U��+y��s���Ap�@Xdt˥�w��:Q~u�Ճ�_.e.K�9�Lb?p�i��}��J}�(|TY$	���Sx����|B$9���LTS�>���z��JyIgn]��*t��*Q�k,��F0�z�`�6��]I<�&-�#M�3ޕ����:
2ut�U�љ��U��Y���T�`/=k4��HE�$X��F ����K)��"��'�v{+v(�M��-�nѪa��O�61h��$�]����\K�%��Y-����ZZ#t����L�'V��`!��
ږ'=y.I�=(����:WPǦ$�\�wڋ\q����s�5gRuG𭶳�Z�Z�%�_�K��pky-)��ϑ0D�ԁK�1e�}�J
�v*��a�5=���s�I���of1iBf�6��?S��\��S~Þ��!#N�sM��{p���ze�x���GA*h��4����<oa;����[�{X:i����s_'Ŋ���X#��I�OI��1ɸX��)RUsaB&F!�ԛ̕e�!���*�,Ē�Չ��@s�Z�ʊ\�͙�Sfv��@�E�	 ������b�}�c��kQ��X�o����-5�!Jat��;.NZaHIK`լ6�$�Q��gʬ4��%�<���كd�A�wT��W~1�Z�đ���H3\=���1w�.��@cEs]���u�~$Y�Jd��o�D�]��fW���G�QG���$D#:�S�ʩ��V�Dmj�4�t]�U���IT�o��Ն$֘tB�.?6j�m�����%o��`�QV׫���M���
Nt�s��r�����P��}�ƕ)j"ooMRv};�e��h�^�K^�Z
s�]��ń��N\�T1ڴ=�� ۑ����W��uv�cb8�]��νr\�.	a�ִ������:�x�Wy�K/e.�u��[�[��
η:J�&����W9�"��#��$_$��?|M��.YÜz+p?���g��/~b��av�Ha�Msm���!�P
�5)��� (-
_�}��H���?��*�b}�a&�)���a���hc�u�L����8�O ���;�&�_J���1�GBZT=Ác���?/a�sC7b h!K�L��D�=� ���Z� ��=��Voꜷ:�i@��#�Q%��pl��}�%S0��N���N� �W�J͜U^�a]J?+B{íQ��SS��`���ɔ���z�H}��kg�McWy�s�c�к��_�������ǲqڄR�^�SrC;���P�@3�f�䣶:/��3��<2ܲ*b��{��)X1E�VmX��ζbk�5`�/�	*ϫګ#lJS)#c���C�{)A�E����\[���]�ڟ5�x�Aoa|��K��_�1��|�/4����^o�vȩ�
��ԍ���s%�-�u��4�j�k;��z�j����~�:<s����PV�f\O_J��9O��]_rv��|4P��j��k$ѵ�}�,��`�S��o��.�ʦ��o�
$	��jl���t�V�E��;��؂�!�W�M�k������E߹g�V�� �ɯ������Z���*��\/�6�kD*(�uV}���QaP��Gv�|���H���_T%��$� �$݆n�L��OK��I\��X8�ÕO/e6W�{E^�ˇ�
q��6�����|^V��"<V�3S[cN��.��������r�MC�A��8����;�=t��1	�Z,���f��(�]�'�;��38?�Ƴ爵9!Jbt8��Vg}#"�>~Nqu40F����������_�/h&�.��r9&�� Gs�b{��*�H���j��qv=.Y܀	#;�����AXN�i�<]�y��ɬ�0��HA�t&[N��QPY$y$�+��}v >�5r4��[̭�8ȉ�W�x�{��#�J�0T>���3�DA-�������Ș�|:u��S
�!�cu�)�a����?�JW�!QJu@�,���=0�`�p���es܊�{Ju�5�+Uc�)VL�$��z���-yuJ�z�=W��\_N�-#�9��:��l��#��D��<�a֛���C�9�v��i����4���\��,i�M�Y��^.��O�jH��A�D�p}��v,P�¹s��]��J���S�ɉ�T�?�X�ݘِ�Ꟑq(ߜmn����{ȗo��~��%8�5iV�$��i �����O�@���8����q�ULÉ5�!�i����N
Dv�d��\���dP�E��֑�L��|�������r����C�D�ma�I��,\ՠyع�
��i��xj�?ft�ܶ�(��k_�a=4lj��j�YEո�f6����)<��:N�ȃ8�*,���'~�������l"��,m���&��ࣜ)r�TQ��=���iP�f_Z�E!+&9�=3��+�$
<&��Q�:�w;�ϾqΘiR�s��}��.�����/��xM��MXheZ����������4���x�Ȼ�E���@2/��{Ʈ����o53��J	d���L�:�z�Y ť�VO��-�(�!G�����h����θHƱH�JJ�U����Ϗb���ܤ��� ��j\���4,� ���RPמ3�q
������Քa,�x���Eύ���aE�B�F���JNL0�	�ej�4Í�Rd2��Þ~�,}�|��� ���/�2�|�i���.M7�H ���U.8Ԣ�q�%e�Zٿ��ڴ��X���Iװ)�������{��	T��-~�h�k����+�����"�A{Pow�׭�x@[
�q;I&gQ�p�Ԋ���ЁzJG.����H-Z���-���:��'�gx�ZOR8�� ����j �`%��B��6g��\V��$���R7/g�Lc�"P_�&�J�q���f��8����E� K�w�/�ؖ��&
*�����_�4f�I�+��+ �Z�i�u�u>�B֐W!x��2�s��~�|�
�J��qx���i��V���˖��ἁ�4C�X�A��)�!>�R����h�����.e��2��F�w���[G��j�������j��{���Χ��5�@�G���M!��֣�Q?Įp&NB�q����@b4��G���
�/���i6$�F���}�wlHz�?�>�p���T���s"�t5)@E �-ѐ41��wĝf��suY�����c/F��̵��|ml�߃�S��:��gl�kH��)��Tm؎L�u�ԂrZ���u%av���n�/v���*����$bR����������e%75�u&$=^�--�Lq	��� ��Zg���U�����4[��4�D:(ny�A�WO�yԅ3R_�$�>^>�%��8/oj�i�&z*�4�I+�����㖘hr(s����g�#�@�t�܋�-A��/E��X���1��$��������J$�	4�0��VIe2j�aZ%f�%��x�h�M�HR:��ȭ!-�	�uN*���&�JhД���U��"�<F�>~�R�wl�CF;YK:9-�+�ò�������G#b�ւ=�3��.<r1���9���L��G�n r��UK�I|^Z�d�:j�#��u��^�a-)a�C��ُߘR���S,�q�p]��|��a�,	��K[d:$C,Ã��ԉ_�:�c�c���^B��Y3�F`k����M�hi��'~�V8$�e+D���}=k`�P!)H;Ս��U��g�Q�o���'������G��/Cæh6��rď��������Ί�pp(^bP,�ʢ\�^�r��)E@�y�V1 @��@q�N?��/f������/�Ŝ�C;�.�����<4�.�F�cw�~jSZ�O�A���>v���M�3�$�x��uZ��I5�ܟ�t��"�j��R7{7(��>�P�5
�L�C�Wf6Xv����P��HJP5�ʮ?g0r��<�S'�n�C�l�iti�=HkKЪ���P;j��f�k�W9� ���,�*�u�(7�p�ɡw�7�G}z�ڐ�@J��R��N;.*�V�[�=���;E�9�&m.�N;���H����g�����w?XA�V���!��@�2��;��Ϻm�y8��.�*PZ+����%Pr���Uʽ!�@��K��, �A�v��8��0�a�[%��R��6=�cSL
��s��4��3I�E���Ӫ�O(8/P���{8;�:�u[����Rh�ͷ����/��h�/��i`����A�Cc<0?'0n״���)x1}� HB� ]��L�R����y�X����~~�F��&8�f�n��u���F���QݩC}�bK�!'U���	Nt�Ѩ��m�aЩ#G��(�w�X���]�Ȉ�b�4?(��E�N�!k(g��Ű:
x��Xz�Y�&&ц}o�����P����ct��\�2�6_�m2�Ezm�H�s4]��C���~����ÞJ^�a��d���T;U0:N���E�+����!��	u� b�yN3ڛ�S2=#�-��9�|��r��h�M�R]�Bb���q���8�]YC�鐝t�QA;%
����7��b�n���k�I�p�7{0�3k��D6��!��f�@-A���)�#�1^�q5%Ĩ�Fώ܌��������?�;,���_��������D�����XdvZ�G���l�u���y�!"A�8fu�7}y�����Tɭ��(b��q�|�{�]������q|\��/&~r�O�4�"qf{)�j�=�e��_�G�0f��4&[�^�u=��\�[���Ck��.)Vj1H���zu��I��k�{��v�1f�O�M�,���:=Ķ�ݒ����SK� ��»�x��>�����v�N��%�h-w޿_"i��?��BlA����3H����6�p�Z�О�"�X��t��#|(+��HV�@����@�j�X-�	��	&��B��xnـ��f:H:�\U$�����Yli���������*g����'�t�](�o.n�Gs���%v+ς���ܠovq=���1���B1�P��ꣁ������z��zQ9����?�ٜ�*�h��'')�Vp�� ��%U|�:�u�Z��x����J��騸I�z�-=�
Ӊ�[��=%)8N���R,��xȹ���(�V85
���[8��a��J9.�}ئ��]v��t���A��Y;h�3��O����PL:�<�s���	)�pj��/�r���s�{FÑwA�\�V-G�(�ԣ�kT�9Vfi%'���>��6�+�VY���YHXiB���������](��R��?2�T{ź�h���ϵ]�봹�S� '�ļ	�w�ʮk)��L����:�,{B�¿LY�pA/(�To
���N���޴K������(M^��7,�<�"%gﯪ�ɦ)j3�v+���*w��Z:Q4�8�6��EF��/���/x�?��E�,ŉ�Ի`�.)Џ�D4`1C��Y�9&�b�7�)�5��L]�Ϙ�ʊ�Q��]/ch�;�{�� s�Y�z��o�$���I6h�"F��e�xt�н������%�^Һ�ʙ�$ ��!�i�Ʋ�Y�B2�[���XI2z�uXAL��;	}��qp~s�k�� �hH���qZ��ڏ����q�L�1���t����:@б�"g.�׬Vr��.w�$��J �["v�f|K_���K�XWv'�/�F>X�W+	ٞ��E�n
�x���`��WH���gO�,��+�{v�3�� ͲN��]��0.�Q-eQ�N`��๝��p�a�H�yMv���B=�F�q�T��|i����X�<^��8�H7���s�|1�B׊��Qk�OI��t�/���^��ϭ14�e��!93\���(F��t�qjj!o�R�{�u~�4���������\&��죦ϛ+�����뜜�Dx������4
�;4x���ɻ�ߙ��)	ZD��R�G�a�g�5�	Ur��:g�H��3V!̤����8H�����8AuoYJ�l�(�&o%)U�2�aV�L�K9c���}�MݯJX��7Й�y!I|�9��c��^/=�=�Q{��������'5v��'��9���3
א�|��y�����F�~{ϯȸ}S`�����<J�p���A�&���,+>��\����%�LQ��g�J^�����.Ĩ�,�Ecd[��>z5��O�CUj^_��8����l�ҿJ��&&ηS��\P��S2���\k��BH��Dh}�mXڶiB�xޒ��������XOT����i�If��'~)>�����0����ڎ�;e�o�ӡ.;D�x3/��ưH�!3:���?���t�1 �$P�:5�n�gKeZ���vn�\n����,��(���_s�y�.>$19ɾ�G,���K_'������� |�$I�30|R��c5F�ɨd�k��4�pj��`�||��=�|��H�x:7cD��kw�q�ə�yHc/Fբ�]0���Bg+h�|9+��c' 3��<·_��SW��z���7pm�&��XV׊�'�
��N�tΧ��CH��^��2��H�����YJs�=Ϝ��A�|�ޥ��x((�����4أ���g��{_��� f��SZQd��'>#�Y�>��J-�䪪y"�I�8t��Q�zf���t��R&N�2��r��k�򫂭�
ҳ�ۺ�i��p&� ��k�;6)�Hu��(��,t�����ݪA�-`E��x�1���o.HI��M@�6�Y���8��<ܚ����[:��#�������j��kK:��b��2@"!�=�瘩�l!�fm��+M�vjV�p-����hLW�U�#�үG���$�岕�KF+���	q(��}��I��(l��)���3u�����5f���EwQ/��-��q&��.���}�»�ֱ�J�T;���x�g�d�F-�����K&��Ծo�k=)ؼBᄜh��C����zƒ�G��~��
Z_x8�B�a��H�<��~l�!d�6���㭆�m��K��Z���(]���������x28a=� �	]���[ү���<�'����5�6��o��~N���ҧ��������K�SJ)�YC=�D�x��q��+�\�ވ�����Z�*��N~5c+c|O�\�G<�=�UŇ��p��
T��9f��s��B�&n%��;��io9~��E�R��LDV��$j�=�Cb�zC��8e����7��<X��m`ޗ@����I ���������5�R��@	��)�|")�i��ѷv��͋�,�w���'ﾤ^��^J"䮍7��_�?y�D�Vʗ���������j4a��h<r75|v[����1�L�,
?�u�?�GH��V�\T���8mVxT��1���]���+�bK��?�x*u��~�pA�N����X}���u���ֈ8���*l˖�M����SƢ�AV#�H���U��yq�tYRA&�8�@��<�,�C_`o�N��D��I�]��C�<�i�u�nT�Q{���ME���9'����p�,k;�)Ն ��\�>���$�4%|��i}��Ѹ�Q)�~鶼|�?/]�z�?��#D��]Cw��F9�xS��B��Cs�.F�2�w�~f.*�ë���I��}�=�����ejK��Y�X��Y�����I��I)p����{gnb#�,.�żo����F�_b"���X��ߺ:Z8zu/�9����q���[��]8����S��������`��R�>�w�'s ��k�����[~�f/4�x�jf4ގFόL8���0����+k�� �-�v�2j���8:�27�zz^���'�}���;p�ޟ�K9��'	���;���3�<}�S5CH�4�GX4$�oi���iK3�`LFA�ͳ��yd����n3$yF���
�$��?������Y������o|o�5�dݚ@iۍ�IX��sV��y�֦����^��%�-���K�w��\T߽6�U��2��+�U���'2;��1ĵ8D��)j(h�I�A�o����-�����Ϧ��^e���RJ/�MyG#K@�Ś�Y�]�
NҠ)H�!������g	MI��_
�*gpZANT�� KiK��ڐ���8C6l֒��ĺ����箹�?	oA�_�ѓ>{lSɧ��4���ȷT��&��.qv)VnK�q\"���y�
:^����*ݹ���<��/�IdW�����[Æ����R�%�~�Ai�v����H��p�_�z_4�WsN�o�Ǝzސ���G�G]�Z\��>|~[Ҡ������DĆ|@ߕz9#D���潳-�	�|]X�+�����Y ϱ`9�v`��\秷J�*!�����?k�E$S��p7#i�����W�<�jHރE�,ukF��)�����/&���\��	2��{:����ޡ���J���2�fb��n~T,�{�L�����$�{��'�EC�Wj���5'����������<� ��2
����Ί��[!�ڬ�18��N����Y��}#����R7�w�nG�HOc|�&�8����������=���WD���Z�\�9��c8a�@����
���IY��p(�7^i���uB�9n�:�)R����qx�o6;�o�v���05�2��~>����3O%�iyz�
G�Y+�c��iv��q)��o�
QS�)S�LcI��!�G�#��Ѝ��&­K���ʪ_��Եy����ԏh���yu���_i���<-y`��(�&����f�=<�5��q$,�Q���s3�
�ײ�����:~/]sA�F摾�=����צ�`�K����^Y?��m@9!ߚW^�7�όȖ�?�t�_�b�]y��`���+��9��Ӡ���+�P�� hA��|P���{"D��i���H�QT�\��3���hU�����S���1 �-%��88��g�O�"�Bޕ��?��Hw���P.��%��Oê�R��w�I4$��yʼ�]���?���CU�q@ !���SH����х%����zR�n��V!��凛����R��1�����̝ќ�m�{2� �=�f�|k��t��@7������}n���`v�·��}���,[,�H�w���X��}��U��^���Y�g6i��#*�B�rt۫δ��c0�x��O�n�Gᅤ/I���M|�֤B�n균E��/����٢ ����f�.z',)�[!��r�OH�
}�>n����y�0��5Tw_���$�^"�=qK����.�ڛ�����	�2J�ό�{Jeu6e!?�ŋ�Kх�w��Q�|�9�7z�7��&A�L��x�c�yv�@�T��Z}�(��旰`$�@5;�f���QԿ��fڐB���Sċ9�W�{�q����ؠ��/R%�)ὶJJڜ�cT�t�dq�s^�x���Kpf/T���a�m��� �;��0X�C���u}	�R8�מ/�dgH���B���Bp=��wIa�_In�~�cTX
�td݊�9��Q�E
������3B����CHr��ER�=Ū�sۈ߳S��J "��г����#�h>ku�2tf�g���ƅ������_�o4�iJ�WV��86�wM]�8���н�4��LVm�?�?h�˲� ��h(l������3�3���s�p����M�_��>r�ۀW�믊^!�����+#ї���HSۼ�Һ4�a�$aM���h�f���]���V JF�b!�b#��D/D~e&o"���*��9�/1�Z��������n�tG���"o���=B?!�ƻ4e���ᆭyM���N(�/g�-���r��ķ�ɐ�n�7�p����?��ֻfΞ��D
�d~!V���h�&�Z�ƞ�F���v#����F��}Hz�H�1���*��Dg��ϥ���3h���A*�f8����!L��F��E�c-��v|X
~Ծ�nݣ����~��h��X�k~;���L0hT���k>�n���N�<�>@����)x荠�7O����͝�R�S�}���D*�=M����g}���VId5�rT�
�E�y$!1@�ǉ*�,%G�p�蘏t8l]���$˓�T VF;#w!����\=���;�t��u�6�:ř�W水�b���Ϡ��WO��D/�eכ�^�3��Ө�R���b^����A��+�b�Y0�Cr�qo�r�,ڳdঙ^�Lkb��M���Ǘ���s�U�3+��*�gy��ݞ��5N�?�b� ��i�����ō`�����D���˅k*e#�˸�I���oS{D�U��THJ�)���	�}M�xA?&.�yv"og���4�8>R�1߼N(�x<����h�9�)�unE\�;cJ�2�N�#����;(��qc�H����my��4`�S�t}BS��G��y��K,No�m��\78@�1#E�Vp�R�h��R��͜� z�s:����)�B`9�����*�����F�i��3��xO�����*��m����M�~58`Ґ �b?��M����y��hP��y\Y]�4oH��懶��
i�K�!��9�_�{�kz��4&�r8-������E�dHp#t���(U�a;;���%�˟I=^�����/z���	�����[�~�]�6
����_ ���Ȁ��7! pd<������:���@7m���	0Ra>e߉�"n#��bf�A[���짳Z}�<��ĉ�B��ͦ�� �ܒ�GH�%�h�|tě8���g�#T���U!L����6}�5�/��?����~��������|�}J=�~�]�)d@8�i8n;C�X��q��]��?}`��vY��P��^�)�N ,hE����(
Ƕm۶m۶m۶m۶=sǶ���t�a']I���DP�����$LA��`�Ŝ矤cYw��yu�O���q�#s����67\�7��;}՝v�;�K`Ι}�{��
<b������4)��NA�x���V=Z
�o��_SM��ZV��vx��b��މ�N^���<�[NY��|���A��,ن'�Z�B7��V��b
�y��O/1P�[��x��O^��UiӌF���`h`��B�#~(֠�2҂8��6���H�{-�L����X	`�^{�����bH���1�z���MR'�k|8��M�ҟ,�O�~w�-x�wQ;��Q�աI�5�H��$�x�P��mw�n�l9��8�����5"�w�!CBw��Ғ���m��dy� P*�ͤ��E˼\����M�_������(�T�}����"��T��L��o���e�P���K�`� J/$훘mse B��#�{��%�\��iE�ho"Q+�c&�u�<gQ�{��uO���t1gͳ2%),��룻w3��'h^KK�%�R'����[ :��
���1S�H��� Q�$s5}�K��(f�A�Dx�{J���A�4����19�V�Gp�G:
��DDY]$Y�j#����(\a��|�[Ѓ�n~�Dd�z='�˨��M�0xn<-Yn��,�Qd��Ҽ�P>.�я��'�,��_�� 5Ma��Ux��t�������*gZ� )|F,F��팻�Mz*�	^HB?y2�
��
���ӭ{E�d��aa3�E���z��㔏�U�.����3{�P��dOjbZ&��.�b�w
}sN�O�P��\军̨���;�+��'�����]"T�
���EO$<@ϴe��ۂǚf��b=��:i�;���fӪ��.�e��|�{͌�-	��$h	����+�'>zJd#�n���Vz;��L9��Y�.���S�:#
h�U3i�{0�g�ˬ ?b�U�A@�	�����ׂd!���v=/��`���Eov6v�N-�O(0m�`*|h���Ν��q_P�ܙ-YͰdY;$��Ok���g�fU�PK���0����4	ֱ�~�~"p5���xQ��D�U�}�p�<������2oW�T�y�M�.��5Ӝ� T�4�#�<�E�2�J�e�Q��M����i%�J��^�V�5Ŝ�ݥ���+�MK)x��Z+f��z�l�����B�9q}�i���L��ofz"x|z���6���f�Q%.�X�m�� >���>1�+����v?��J�k�t��񤥑�w���V�Vˡ�3��1W�>��.��KF ���G��>��U��w�y5���m'��R�jI�(�u�Ta�/��W%=�����d�_��Et�evRge�d�2��;h�3�2�2��DZ��f���5Y�'1X��n(�gR=$��^��5�6�?��,��+$�KR���J�\���zf���xWV��a���e]�?�?>�7�R�\��P0b����tdNg�)�w��I�VS&�n�h�F"�ȡ��K�XJ���b@���,mp�b�AKr:�4�]�A�P.:��L^���Dݠ���A���n/�O�y>>�`�����A��3T�Z��)Ӿ�\��o��"�}�G� ��#�?*̠I;݊ȅs�G��,��T���;�|��/$�"sg[�p�CyxT�1c��QK�Ʀ�.�q��rvc�����N/Bۉ������i}����ks�n�^�Mi�
f�c�3[�Ҹ_�$!��E����_����?��й1�Wl�3�B�^���	�K��VL؁S\�7