��2���
ˏ��Hy[Um�����v�b�5�s*�l�"W�]��h�nGF�����[)L�e�S(sy\�Ω��I>î)�GP�/y�j��3��nT��[�N�n*x�D��v���i�ݡHZ����9�ꨗI�*�mY�m`�gr�,P]�W�Q����������,Gbb�DL��DJ*N���eI�H_sZ�t�-vB-�[�V�����9�u��`Gg'Ҧ���:U��g?r���R?�\�c�����#����.�!�I�r׾�i��o_\���Ge�E�NWs��s�������^BxGkmč���d��NE�O9��&X_z��0sR�����7MS�/�3e:>�jb��o������9%D�kK{��=vvVh�"����_�"@�դ��D��'5S'���I�q�I�C>bC��ʼ.�ik�&U֚[�o��hQ��i�g�BQ��Y�a���5ݑ����՝���s.C�A����m��	nY5_��uc�K��oz�_���qIW�ޣ����W����x��?�{c�uߔH���<x/b5�Z����������벖�
"�ic+�	

�
�RB��k8�[�6���i̭<,��ܖ�0�9ví�V�\6�]����>Sys7kg'wWg'px)�mP$A�Lo�Ez��1������KF'���E����m5��E����k%���������*�|��i���.~��@��?�����1�_���!��\�W�����������_���o(�����Í�������Ԕ�'�]�� �)��o���7�߾�5���ܚ�r?�X�����C����Up/�O�ͭ���g�_�����7�o8  3�A�~���'i -������z�I���4� ����Ȓ@��Y����������J4��7�Ńn/'A%��ܟ]J�-�����8��?�'�cW�N9|;�(�e�爇Ê�z�|����,�a~�����E�?��%:�9�i�i�d�	��rs4wpൂ^�xG���S��Td?��Kҿt�.�,���U�jyWc��������|�^~Y;���s/�[sknͭ�5����?�������k��L���,�OG��"�ŵT��hq����#��@(eg'w7���#Z�a��_1~ܥ�g�u��YŌ{U7(��b`l�~A���:>(ŝʱ��a�s�^do���)��K�;�G������q��ٴ�D���.[�ǽ�	�_];d�>����QW�9F_}�N�_']I�E�A��c���x�8O�]+d�Ԝ�3��5�:1�MP��Q����,Â(�4��/hQ�Q�=_����%5�������xt��z�|��ga�YՊA#݊~-��}	�9�{�Y���v}oSA��
+m2���i�o��~�� ��7��V�±���c[�
Ƕ�'�m�38�2ql+�±�Јc[�9�m�q�
D8��pl+x��S������cO�ǞB�7{
���)L��SX�cO�Ǟ� �=E{
�p�)8��S����S��߇'���@0�Ҟ!�J{
�ȕ�yV�S _y]B<qx�ᱧ��N�:<�����]h����(��B��&�N<v�w���c�a��J�	b;"���W��� ����N�sO�ƪ�q��	Z���"�H��\��ڼ�5 ���W���0�k�:� �LǺ�MC} �VBmj��&��XJ�<:C3;~�L�uƵI�'�q'�B=���śU���:�2��*�t�+��Pu�>�뎸33a��1U��h^�Ull�l0~�&���;�j8ۺ���X�#A�f8kЀk 5b�����p��?>v�,٦�b���lYc�3��!ԠDe)2"�3$KS1R�(%���vR���2ƏW��,=���}��������=�9��{��y>�AG��I���6�s�>*eK2��qlFk��O
��%̳�&���I���oj���ju�+oO��f�2��I^sg�jR����(8�>9ȧIU�)
B��܉�����T��X�V}浾�
}�ɱ}�>?|�g*�@|�# ��E4��F&G���B#5��>�>�p�]讖�&n�g��RT�ˈzy�k�,\�G�����̼Jv󁽜1Mʄg���p����VL��1�TEG&���bA^��M�yj-4��I�!�ƃt'�{��?qW�mjߏ�~FT1ֵ�����.WU�ϩ�`��$���r�
o��{��	�f���u�C��-�����ß�3���e�Y��m�Lr0|o�z��H�s y�v~�=\��������z��|"�( �W��r��{��=^�Ha��9hŏ�dja��Πw����g�����x�f ( �g�������t��ٛ�������_�u]��u�WDm#$A3����w͓�1OX�k��Y�����6�gh+.���������������