Fg	a*����t��qa)���Jq	��k��wm�0�9Z����g۟IE��i�G����%N}�Pgäu�xۺN��[	�B�ü>Z�c2Z+�
+y"L�״	��_4�C ����:�#r]ǽdwbM����@��	7
��ґA�˓d����T�K� a����칸��S-��s	.�N���P�>4�-Y ra�,.�5�H����G&B�R��NfS)�a�	��]�����|�Dת|u����w��"�̕��e�ȺMVb�Y4k�U��m�h�7_���QK���ȩ7ֲ���Zg�l{ƥڎT�Q����vK�.Z����C��b�_����j}�4�J�9��5�#�]g4<7���H+�i6u$r�kӆ��O�fZ���J3���6&�x���M?u�����Xw=�b��������P�2���J����Qy򮇞sU5j}rK��ٮ��g����f�����vn������2E������b�j�"]->ᐢͲ�Թbq�}m�+< �F�j/'����vK��.�3��k�g�^6��}�V�Sk��w�I>ٿ�LF�S;�"����W�����6�{�L��k��R
�trR0~�n�K��V	�j�B��N�ɼ�O;6t	�qt�ݣ�^ړ5,�ɶ_��*t]�e*Yf�o�9��e͘b-G�z�n@��x[�<t�C��?�b{X �G7I�+��=r�v�_
�H;�:����v�ۑHW.���B��;���a������\{,��+�^��^ �u�Jh̜h�0K���P,����,C�^-���/��8����m�l���Ӻv�^+����=
�{D[��WJ��������Wޝ1���06�[̲��U�6�՛y�4�_���q{�~�A�iZ][�u�M�ؚt�F��:�o�a�^T�W�M��]��$�B=S�u֧��$�aCm9׸�mH:��?V':�?�4�u¯����?p�N�B�}Q��ʸq��n��g�Z^_k�Jm7&��'_��u� ����w�P%�c=Q��OWH덲*����܃_�� c��܂ ��<�!�aY@?��Z�:B0�d��w0�1����ׁ��p�Hg�^�\|�#����Jo����f��{X�`�|K�<w"DA���c���i��l0��E���!������� �@o�����|��/������#�1���Z�ouY,��ҝ�^��ѷ>#/� ��5�ȒO�G�j����u�+��;���w}�@Zw�$�R�xSV}�����W�Q\��l�ڵ�7�l�+���~q�]���b�������'�?kp���g�)�o��9�o�Z��)��M�F3�e0="�5����ڇ��N���'p��`�}eP�,��ncK�OiYW���R"��NG�b:�[��{����N��'x�z�o�I���O)_�1������/I�$(�/��Q
�����;K����M\r�+8�km�{�('8L������{�E^��&��H?VV��ܹ^�Z4�8��+4�z!���J2;��+��,[$��K>��ɉN�=!Ƶ35^�%B�G��[ϛ;}]����#H�Y]�X���v��}1��G�M˱�bƴ�}I�%@��yo����D�"�z�s�nU߮��k��#�	��/n���J��b��� _D�� Z�y��Q�Y�(�E5��՞M�W�w��b�d�~)�=տ������N���2 Z���,GD^\�R���ϻbW�D�D�	-���ϲG%��{-c��"f�r����X����)��?p�e�����HYm�c��K�L�;�-��ͯ�z�Z����?�XIe;��4E�=	��x�\��vʲ�]n&khoF�	�Qm9^f��8�=|�́҃�Q�?�['�#�䇞ʿ���fH�t�o(66�L�SLE?������U�w�K�v]�~�_p�k�՚p�ҟ�"�%�6J8n�3S�o׿���y���������*_l����� ��𛭆;t�ܷ&R>Ib��.{��?c���#��q��UOU<+gɟ�T�mt�;f�kc���j�q��X���~��k]"XT������:[?��gx��ץ�\5�?ӆ�<w(�%��w_IDI����W��ϻ�W���>�xl��ݴ��e��D�t�x&�K��E?ppVA���Vˇ�c$܊��[�����?��^r�5"fi:w6m@�N7]ζ��Z�<��x�>��,-B�u���|�ѡ#�����-82'{�2����i�=�{<���"���X���e_T;8�>ƴ�����G�e	�%f��?5)c�y�	��n���d=5�zt{�����t.�\�J�֛2P�>�	#5e�t�jб�0؈"5��x��U���+f�a�'�l8w��j�-