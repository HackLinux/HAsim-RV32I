�3
�EmH�1��̛���m��|�C�E���ڕvj�ɲ;��_E��uem���������ę�Ǟ�Ɵ�Ř�̙�Ϟ�Ο�M���f��-GW���ycB��S}��n����5�)�ҫ8B7��y=������lG���ˆS�2�W�*�C�0��)�iE��Ӱ$s[��v�������u
�u��\�?���������>$Z�Gߧ�����#4��*�#-���.���������"�9�=$�{o˩*���?O`���"�t��b	4���w�,�ФVe38嶺ۘ��r�����HA�;)īl$	4%���%t!L�T�D�=�d� �Wi�h��
�mAxA� q��� �1��w�GȀkg�"$�Sh�>�s��]��y	�d�h~E��nǯu��9��'|�AvéV�@����q�8�uʠ�j�Ifi�:�c&�Aڋ�\���f��ASצ���"��"T+-�lv��1��ei$��S_�δ��kg����3�_xձ�8ǴY�5l���c.���?���	@����t��p��W.,捂�s�g����UY����O�����BE�S��RX�ɑ��NJ��g�v}��~I��;�#�b�����U7S���d�i�
R6|�ɒ��J
�f#��~����N@�B��H@z�$���<����E�������N�wߤ%�#r,�#Izk���tv�g�+*��#��"���4���(_��%|��T��#���fᲢ��=�DF�w5��Q��.Ӈ��(*"�p�I����e;A�x����i1������d1�	8�u�Cw6��D�c���.��lGk-��V����'olïĆ$&���Gl4�	*�󦰅��4^�ϗw�J��K��d���
v�"�#CA�+D��$�=�N�Ď*db��8I^.� �n�Q��TP�jF"O�Y��N](�D���p��b鸛��"
��ͬPկ$_������z�y��x3@���W��iR�������SG��m����(u�����
S1�x�q�%��A�>xd��%?�ox#�r��Ǘ���m$8�u��A@�,������	��Or�~佾t�q���ŋJq}hbs#�rߞ�K�ek���H��(.�LG(-���F��m@j-�PY�A�3r�w�
����Ť����X�u�`�d��^���[7�ŧ�:����#jd�~��ʍ$Ũ�ǭ��vp���݊�@�~Qdq	�s���N�m�c��7UW��n�y�Ue"��7�6����vy"(
h:|@�B��0���z֒}�;�cJ�~��%e?#['��l�O�ò>�Z*�d�~�_Ն��k������9���gc�Vc�6��g���Ტd>9�50���鈌e���_x%����4�g��0���{7���+,����b6�Jq��u�HqD��lG��в��ᵁ�S1Gx�6�� aVY�����r��ע�������&A��<��a�7^����6�U��H��$)��,"El�����(n�$-�B�y~�lG��UN�e���
S1��r�H��]x%�����)a���i��&d�ņ淄e7?�Mp�d��c��vY�ȖV"��2��Q�Ifl(8XB����;&�fŐ��@{b��|��zP3 ��q�{x�1�v{��A�������K��k�I��=(�J�8H�&�abfe���wY���6���~nĮ��;�t_�ϗ�����H��;.�L��I���.��b�U�]yҰ[�������?���p �*�~~�hy�q����P���k�=�
�tV"dv�Sh�AW��x[%�ׄ���G��W%�Pnw֯��ϯ[��$���;p��I�vA�TI�bM�]����@z(��y�
�>�.^�#]o>��K��4���u]��}n�[V��Vq��2I���Դ���"Ə�Q�2;����J~�@,�;�P8BuY�.l���Z��Q�[�-��R׀���#B�,,d�_�Z\�Q ���-�~��P?��72�����?g��/��x�2��wp@��d�8���>�-�qM%��)�x,=��/mH'����ì����E��1�-��m��/ �v����/[Ga�����`��|l�����_�� Yh��
4 Z_�sY+�&�o��QP�W_�o轵ā�z~������S�IU)i_�2Gnld<�L,�p�(jp/��_<�r��&,|֮��M��[>����Wx������ 8�+>�	½��D��]�Ŏr�[�l����9�v9E�MP�����<�P��EtVA�D�� 4]�]z�H�߳�����; ��E#������%#`���	87.�:#��Fa>����X��-ވ�1L�=�MoKW)�ˏԿS�^;U��P�)�{W��c�@c��yʴ�B�`������?͜
cYvl(~��dN�J1W��{���<hf�?G�w+������wD�3��**blY��S��F(�(��S	���0'Šz~�������E8�Wcz@�J^[������:�sn�I�-Ks�QR�`-C҅i^#@�_�n�?���
�	�Ki�G�6��CYs��J���:qsi��I"�KVQ'�w�'�gޝ���n���_�GG��ia�F�Bc@��s�OQcƎ.����>�Ү>�Q��e�����ׄ�sɇ8�(��=�8%����׼�6(Y����ٛmao$�6;'�0�N��[�=�� �1������S������P�+)�1rځZi�*sa��^��<��X�M)�MY��R�q�O1�+ �����._�r�IN4AZ�'}	;nZ���|Y!��������@k�7��gX8 R�6\�$ B�,,dj_��Ga{C��Lo�=4��?�S;�ǯ���8��[�W�|�u:�^����s���;i�6��A�N:�aN�a�Q�W�U�9ב�}��fd��tX��}Ok�����b�7��	��/q��,��8������0��MV�E���RVF]�B.�H=��c�Hֶ�X��:��<j�����b*��}?%�,�_ϱQ1�8�l��ݞ�NWH@n TůV����9�0DWFE.$/�F"n��l�Qi@�i/��(U�_>D��vV���DT��`�K<���h�H,��V�q�G>I=l~�T�J�$�H��s�A�e���ʯg�8�<[�*�z"ǭ��F�v���Q�ʆڭ}bn&�1��ՠ��ڭA���4eb3�Oc� �񢥽Д������,&�&���j�Eb�1ځ�\�%-��mЕl���b�.Z���[b6,yĬ����,��5xw9�o-u������Dl�����Li{r@c C,�]\lV¾S4"��0Z��N]��׍����.U ��ŚjA�8���M�d�\\����������g�[��+��o[�"�nl�g�Lt.q�#�T{�ёi�����!hM����~����憙u'��V?��|)���O�H`{$ɲ	W���q���� ��n�������q`z��T���S��6y!���J�
P��N1���l\�zó:�)ݛ�w�G��N��6����n A�j��ﰳN3{��1����M������bPj�UK���Z�]�BwmWF�æ�Eu<Fq_��a?�7��m�s{]�Hwk��
�J�p�m�	Ĥ��<�ׂ�=��e��_K@8
S|զ��⁍.z�^9�J&���id��>��ݻ���J} j�i$ D�B*��VHDT�z���n�fz
Gh���`��Z���
V�I�)a����!
Fo����\�,у�s?���o(?�Y���o4�Y�_8�Y<�7�J9���Gڙ!Hϻ���(�^_�	5 �~H��ɽ�NV7N0�M�)���~��.A���?�N@��o6�z�~��1I�=ٟ��N�J1�Q�Y�8�8I��Ba�:?�j�@(Ry�JLE�$�
|�Ļ���H>��{-xSD���)�g�MqzI�Q�{����{k)Ŭ���c�a�ѕ�;�2&�jlg��q��;�N���̎�Ofs���$�����Юl�p�\�ܗ�i1�b
�=�Y�
�!�3[��܅%�*�}fQ�.Z� ׋;�@��E.x6/@-Ǘ}���n�����g15�?��0I�*�B
���+8t�g7�h�����B��TN	NRFﻲ@8�>�>�w�C�B��A6��J� �UJ��x����T��r�q4�6��h�_�ԟ�M���7h�,˨C .��s�TNA��<�kk&�N�5�Ɠ����vTuRϺuD:>i�|��C�4����� �!��d��z�'{CS�$�i�`}=R�����_�ve�M7��p��'��ޚ�E�"r%��o��I�����=��q(rg�F�����ܡ��������}:���O�r�1�fH�浳�'V	��A���׊| �!����b����جr�����B�:j��uF�D���\����"