���M�����)I�4�S
R}�C�ɢNW`�M�c������rPsWI���p#e��Nh�����e����n{�2�h3E���ðܐ�q7��J�0	�C1�l,��g�X��6*���W(�ܲ8�n���u���M��/���Uu��T����);e|4����T�Q�������H�c� ��O�f�h[�Cؕl{�SlY��4|SD!G2T�N�e��E��
_��=����ݠ���S���d��p��|���:4D��a�!V���B������`�<s���=�����cm���=� ��D�gB'��K�۲66��4O.�D�����d���3����7<�U��1-1�I�O%Z ����d�8�`*��D�b�#`k=CB���Ni�JB��ѪcF5R��f����)�4�|Y�ZR���R����l;󄦵�����c�����ر�����V�;i#��U�A�*)�OH�QB#S��U� 3� �ڬ�Wbj���Q��dŎ����*��C��� ��V��Z�Q���w"Y�����/A�����i�ӋB`;�]�v���\�5�����@C`"�N��h��dg����F�m�"�M)��s�@��K��^���lN���T�����R=�!���	$�6���}#�����ޓ_�>��������g8�D"�z�6�1�r����3����!"��L����=���������|(Τt#60��H��Yà�s���������|�B���d����o��2��R��C����y9���9ߴo%l������c${#��l�A�d��e���V�Al/���W���~y��j�I����ʢ_g��/�G�(�nY�C;�]G�C�(����x�;(���D�f�]���r�̤���B��嘩�K��N���M�B��p�`���U�]�[��v�-� ���N������@��HBLͤ����hjs:���헦M�È���%��b|��x�lRI��Yr��p.2�(���v�\U�q����S~�H�`V�����z�6Xg���f�����ﲼ�r�b9 k��#Vy��[%"GxD#ެa� �����1%�h䣓��u���'>�a�-���rA���g�P>���֊���4>��p!����D���z��w�e:����Md�~�6JϤ��>���n�e�E��u�li�"������0����dS�d	#�����R{�H|+̤���.������P�D�q��f5a砗���e�g,^A�ױb��!�Y��a_e�7������ȏ���'���ʑ����爻�»�淠��d�Y���L�i������3̤0�m�f .�t���0RxVy���U�4���X���c�����m�t�ᇠ�P���cm�c$���O⒜6�N���q}�+�X$E��~ܒ$� ������kq� F�f���I����?r�����0������S��B�/c�z槉���R��C�!r�}��h&��{�^�7��'4������E�eB�2�������T�#:R�����f҃U�G�i�e��h� \U�B�=}���B�*d�����B5ދ�72�K�V��`M�5}�0�$�4�E�Ob��<�����o�`:�3���i¨�u�dK�O)����I:���<d�17�R~�bF�myD��(�����s���A[�݈��{�����^��D�f6�֬�e1��)AcP�S�/,�r�rS�-��L6d��C����̇�S���_�69������f��,d�ݪD� �c!��w�Cc\t�$�k+�QJ����r�+q�4]g4�B:�l�3��Dgq��3�+	�>�K7�*�Cf��ɧ��,OP����f��v_+�7&e�.��t&ʃѭ�V��Ѣ{鿆?${<%Ԉ��d����dh��C-�QY'1C����`5( ���KV����K5�#u:����g���Ge2�7M�c���e��������ǰv���k\#c�.�O�d 3,���d�䲃ߥ�ѪN���*��9�1ͣ�%��"d���Z�X�O����@E������\�B�|軔��l���<��@䨉Ӽ��Q���y�i���aj-&�I�vX��\*��}���H`�&�r��8�����d�P*�"g:!�Z0�Ϩ�#żb@�?�<�5u}�UV?�b����3�%����A�།ڑộ�Bg�y�3�l>���z��@���ҷ罢���k�E�6�&���mU�.Ag�Bf��:��^�]`��� ��f�Bfj��gxpcw`������vTu��珸k��[ͥ`�a�^wE;ve����#��Ǵ�Č�8�� �����E�2៯���~�c㹙Ń��l��˝��V�K��o���Ԁ�ǅ!E$�#a���"���B=���l%3���1Q3#��������{��*,� ���D�Hab����bb�z�#��)���t%��cZV��Z����ܠ�(�{r�I�s&K�$� qc���k� ���ݑ�B߶��Og�۳�G��i �б����{��H��ۡ�����fP��o���7�0y�Ҵ��ڦ�Wc�J��2��a��{�4$�E ��i����q#N��Ib�hxsG��kd��VgQ�Ā���۷�a_����wI��vu��~��/�D�#X��F�BS���3d0g��I>�E�⦅�r<�炧��R<��h��S;%K���l��=H�H��$���+*�*��x��O�%��#��;�<�w���û�Q-�vu�t���cHV�D]�o���	�b��⣀��C>dV��������d�慦X�e�5������q�E`���&1�Č�8�u���O�=#���Ce�B�\�A�	c�������j��U��`i�b���M&����t`���#Q�cܤ>�ep�BUa�z��:�c��U����]ӵ����8h�4�	 ������7~櫇�[�dD�<�e��-NW�0�%"��X⇹�H�:��#�_�c����$�gA�d����z�m�׵�����d��0%�ڑ�������<��%$J�& ("v���v!�́���ʝ��D���O�c����1Qσ
�c���E�㐭i����!������!$Kt�Gg2hGvC �H:��~rô�&4�r��u�<�S7����kӄ �/ܘ�ɏd��Y��&]��A���a�3�yY�$K���� ݫd����dղ;�@}{��o޲$�<�l	����z/_�K6�¶��<���T:�ԗ����`�'�1a�5��|�)��rO�{j���Q-�m\�|��q��EDQo��i��P�~������"C��Ȯ$�w���A��"#S|Lϥ�0ՂT����O���˷�AX�d���&Eq�G�
q����y���@�����������ۨ����ԚD�簨��c����vX�c���#wf7����,�̘��+�P��I,��c������E&�"�X��*�[	�c��Mw�G��#ev������2|�o�=�sy�ȩu�~i��a+-���(�r@Y�<�NX3c��cfǱ���8�����˪���5�"��O�0Àw��(���K�AC 妿�%ԜB��c�E�B�uM��r�a�����d���2�dN��~�vN�2��̣�"�"�ä֥�� ��5��������3��ĕ������ɊX|i��P\����5K�#�������:�wE ��)�W8bh'ɄX�P��3Ọ;['ѢU��� X�<�T���vU��ݏ���Պ��=��ޟ��`���&Q�2�t��ʬe��A��v������G�}@&f���(�e`��2L�C���d�~Q�! S��z� ���.wF�z����%�f�>H�o�$p��S��H�M&&�Ub�OE��ɩ�!`ETG�{h_\ �E!v���z�"#�Vq�gR���['��V�����l#��K��+��l��S����d�|�|`���A�����SD!'�*�ͨ�e��n�Ž��gd���M:bc�
R��`�0$���cVzP�ʙ����6%�g!�U��?p�����d7BE�࿳�I�5��t���S�7��Ox}x�Z 0�z皘/B|swJ΂_�:�ȔM�N��UF��� H�z��E�m6��J�0��M���B ���@�A7A��O�~퇟���ɝ��t�@0#X��۽��pg��GS�*╼�l�.�J��뤛�I7O����e�+��Mx��Y?��tMsE6t����Y����P?����Q�Yz��U��.)¢� �(���6ds">����C��k�<ԅSX�T�#�c�oJSj���؁ՓzĘF!WH�ʨ��mx�����Yч�%a��՚#	�A��t����e�����,u���8�����A������<6��x�H�F����4odTm��|��qP��Y�t+��F�� ��xODC��uY�MC��U����xu���ޒ�t� ��:Z:�/��s'i�j�bvÚL���9������������e\����w�PO��1��2�ed��e��`�n��dc�� A����?�m����bA����^�ł`�0D�"6�n�����C��(Ʌ"d#���P���e&#"#�BE�࿳�����ON�t}������0�Ϩ��<�L����e�!*�IȤ��T���K�;3�h��������F��/b!)��ɐ�w�����1�i
���:��`�!5��"g;�k��e���!��%V|�Uq`AϷ��Q�`�_��RVe�7eAoE&�/����%~��U�Ӣ��ΔL����%���&�7BE�࿳�����ONӴ}��^���ȩq��� �L�e ��H��_��$(��(bhg+��W&FA��d�:�������Pe ����N��{��F�f�do���<g8򾎊��J�&���Mx{��f9��F�c�/��#���y�$�ba��;�r���"���d�VB'�/�<��d�}�T�������&�%]楝��F�BE��3�s��(���d�4SgQ`���]�b�G���7&��E ��)D����S8���_&6�r�O�e��c�p��R�Ty��*��5��ԓ�9� ԣ�����ŋ�f0�c�L����H�/_��+����#���o�����ʲ�Wb�����"샳|�S��<�Q�r�g���d)"%��.ED�Ḳ�:t����HD!G2Tf
P�/�{c(��(5��E�����RP9����t�����u��'�ẅ��@�
�b!)�����w����H�ZT��6�B��M�D� ���`*�  |�/�X��O��Ȱ�v�U��B#��r���D����xN���4�2�������#�v3���	��g�d"%by2�č��y3�dq6�Src���q(����H6��"�)�}u���b�0����'>�Ƙdǧ\RU�:ؑt."���u�/C��cgW�<��l�D&�����g�bb����f��u��s��c&c�cO��� �c��c-�0�������0���c�zP��>��g�dN����9��,�����Obc������펬�G"/>���@��1��v1��qU��{႞)4yuqL�d�S�#��2�b0�h�P���<Z PA7�rP��.}�
R�0���gA��~����89����C�t�m	feȼF��O�D��v�ؼǡ%�!#Cdb������t��mLUn�i�0���ǭ/�� �c����eo�Wg6�y�Tۅ֞�O��bE�L�����g���ϥ��B��rJ��S�� A
����61�EN��4���*��;�~P%H��XȣL̄��Y�Wd��D"4�E������ ������Sەq�@�@��2�*�\��$��m����T��U���(�^��c=��MW���%���+t�Vg�1������ ��}e����c�먠��Q��i���˖�ϕ$W2ëS���b/��K����s�A�U����x��c��d4��4�!.�v^�9��7Eb9ȣ,��������(Ũ�c���벟�ѐ&�eEMZ�	Gg�i���+���ֻ��9Kf�)�x�7D7�͝�N.�oX���ߩ�/�$"�u��R����%���J�������i{��Ō�$,L��T�q��ӹe��	x��糭ズb����Q�b_�Qb�Sø�D9�5x�ʜ�O)�h%��������Ѱ��iB�����ax� 4V�q��@����.J����K��3��,��:�W$O��YϢK��C��!����:�ᶥ�©�&%���+�'������{"2#����O�b`C�M��Ҏc��6�a�����2�e���B��-�L_珁�"^�)�y�Ǆ����u�S��t@"����뢟�U�hQ局��E:��+�~������~��TM��Έ腱��7���^�#2�t�顐�Zr�������S:�EW�\��nч��nL��������½�m��������`7)�Nu��X��]ϊ���hV���d��b�Sc��4�̗h��g:a�����b0��!��oK��C��|n8c����Uԏ���?��l�%����r=��$P��o�d���%\�u��e7�r��b3�~�ę���6��-�� �����#&�������j���A������v���&I�$U��Ս��(��_�Q��Sc��d��%���ɓ��d�⅗�Ju�|��Zẵ�|�mf[�u�w��n�F�G�d�G� SM���O��Ԏ�m���X���D�d��b�����D	ϭr�z���$堲���Ń���DZZ�|��e�g����x�L����FJ�N��4�Ϣ?����D5�E��B��cQeMT´�Ci�dy�Fgqݤ��&����) ��J��H��v*�΃B��KY�ļ����"�d#�E��"<�÷�$��eW㘊�KΥ��t����Ҽllb���%eiZ��8Ct�b/5f��,��=Bu�Y���c��$��EΪs�{���(���^��Yᕇ�j������ JblL��r΅.�^�Vc���3�倰���r�p�PeJc��9���<�C��$:�ű�"7�sy�4�駁����7灜�'"$����'b�eH]�yv%������r���
��bGg���Q�$Bc����TR�HΥR��\ȣX�D�鍝耀�)��0��ܲ���'�e�� ��nx]�y�,��@�rH�Vr%�ܜ3Y�P��冰�����4��>���餷#��d��r�R��K�����d'�e�	 ��BËc���$�>�c*��	��]Gg��;���Q刌�U�cW�D���;�{᳛�0)�e���B�����cN!#�P�K����Ic�G����M����Ѳ�e#N�
Cd8��?������u�5��D}�ȴ���j�b_�`dC�� ������
W��en�*�:�����en}t! X���Z��k�d����L�s�s��삼߀���^
r;f�������龕��7�b"���H&5�}�g�}���Ƭ�g�}�g�}�����5�骥��ﱇ�>�~V�)Cd)�% ���k�D2�G������#���&4��p�i����rLD����@���	��KQ�������-r�PL�嶼�H��,�Ŷ��M�j�p法��:i�eF�4R��k�!	3�q����ժ��X��q����6/��x�^P⾋b����杇������?��Z 2ⴔ���k��m FDiM垭  S��܏��{��cN�f'U&T��p�z�Ꮔ�b=`���@�$^�%E����S��v�G�B4gqǃ��~ c�fV\��Vp�Xh�,�sm�p�%G�k��eB��E0�z�_�mQ�8�b��$B�ť��qS#T�$�9EB �����#`S�"Fɽ���ej����4��p���錼䁱��������/�*_�g���[��!��SSú�$i�e^�1������hj��U��>�Io�lD�?c��TlD��fɖ��
���w��y��W㣊�G����s�Y��9�bQS#ZɤN΍�okC������+I �!j���o�)�*}k<����j�m�"N�����)�e(��A��z�Jm���U���ܰZhc���9݅�:��z��\V&�	�������{dj-�Dz$�>�j�F{�=�����n���ۡ����o BU��C��Z��$�Y�z2��	l6�p|.*��S[m<�A7�g��s-~�
�
{��Q}�P��Zl0j�<Õ!�˟|�{I����˖{�S�a| j4�Fu���s���j+�T� $��D���`�~�E�$�I|�(|)���Ag�#�e������%KQ�E�<�%���.\:*��a�`�������y�����6���`z!�
��隈���e�b��������6��Q�Eݓ۝��B�����|)���]�z(G!�{�<j�	� ���g�g�5z����� �p���J��[-c$�{�	�����|?�R} km����>�֛`�\!�=�%P{� �Q����C��ە�B�����P#�W^$��E��S�%cd7��<�~C��tz��	��Z%�h�(`"�f�6�s����jl;���D��g%	#��g/�@���u^=���P�C���2�"{��P���U�"�r�1]5���5��7����l;*ė��&��dj&l��$�+����?�^&F��Ý��/�ٛ�W���R�rC�2A��;���}���>�y�%���f�}����BV�m�d��X���#���_�����G�k�;r[&
ȝ^���F*0�g�.ad:�����E?S�u|j9�z����Z �Ħ��\�q�������|j�c5���3�"`��6^a�oz:l'j#�2j�Q�	�$}�b�jL|�����;zF"�}{6-cd�&�7z:l���&�u���$�!z1l�h4���n�!�+|*��@�i�v�{6�w�\����L{��Ȗ�@_,�%	C��%z-�t�o�z>� �u|b�)�uT��caC�cb�7�{��@�hڄ�
�'�=���4���`�Ë����J}H.�4z.l*�	�	�q����ݻ -�PBx����"k)m!��v�r��j��$�w�oۤ*�%�֚.���g
�	cچ���Ё
��x����Ī�՝&���=��k���Z��`�Z����a�3|n�'���qf�z,�կ�����(�*��Dbh�`�4!���B�l7Ǜ؜��@��" v�X������c��2D��>��#���r�LO� x��݊�~���r�\
j#��+�������E�n�y�uz4��e�c�}�J�V����D#�������!�+���t@�(���Ɯf� �?�q��t�Z{W$�I�a�������\j����ڦ�����@�b�,{.�k�`r\\*
ġ�Q���m���`���$�
�<|�����'Ũ	�2��"de�i��^�J��x�$��~t"�	�5����t2<Q��P�Z0����[�n{ ���9���*���� ����$�:�c'���f�T��TMR�I�yz�����c��t�X�ͥ#���%�&� � ���}r%���`�<�.���f����'����9k.m<����^�l�B|>j�[u��ǝ��H"�0t��$ڧc�?{%�6����Ձ�U�P�^&������k���C������W�l�;Z��N}�lef'�M2�\"*��C�� �E�r�k� ��!+��ǝǥ^�B�N�]cf@��!C��E���-��Bq��ĝ���u[c�@2E�ữ���o���;yv`'qk�O_�E[�Sj����a�t�g��� � �Z$��4�e������4���-����j.:A� �:}��9,��!ʧ�k�c{-t4��>����b�Z��e{�t�4Ɲ�����A�2��Qz9����#}$+��k�|j=�&g�oΚ&�(7+�	�!��\���d�E�k��Ǥ��5C��*#��	�t�%���^���Izl�5�Ao� ��ó���+ۦ�{$���U��#�M�B��"x$�#�'��dD6���8�:���R���2C��\�4�j���Z���R����������]�r&�D{\�q�Ý,������R��[f�]��g=o Z$̡����+*�����]�������	X������4J
s�kh'[#����L�E�Z�3��D�*�b�b��"*(򙄜Sz,.�d��`�"}
su��䖂��6�Gd�C�����3����U�G@��O6c���l�;��f�${u'%�����L��㒔�4����J�-��������g���T���-��杼-��[��Z���u�7��^��6������E���Efܝ��2�[��ZH��g�N\NM�j���C�0��d Z,�F���na]I7_.�hg1��E�>���3HZ$,��\a&\"*�&MBZl��W��h�-��I����hg[c��V�D�;��T����y:i&\"�w�b��ci�@C���_!�\�7f͢�a�-��Z��\��7����$�s'�N\B���6�RZ����� �r�s&�&�b�tR�������9��Sz���:��'T��������Ɯt�u b@��Ci����
S]!���\�:� Z<��S����n�[-��%��0�u����6�d�^���<�f1�n��[�u-��j���%�R&��\�(8Zt �B}P����n�����/�=��M�Z������d�A${\0}9�n��+)�#�[�D�b�G�<��n��[N�q�t`�b}���P�?��r���Ԛ��t���������Gq���W��m&Qd[We���.΁���	�������sJ�������We��iy�D��jR��wi![���f�P�]H�R��AS"�u��ɳ�E#Y|n���m��,�P䜈u��'�r�,��-I��lqf����!����X�H�߮�T;�+���J��!n��rM9�^�� }V(W%�7�@�b8��s9�Uv�a_���魼�h:(qq���'z��!&5,;����T�s�3.���,0�"��:����S`%;W���~��P�h��0����Ļ��F��j�f�7*+���^W1�1�
�Ⴙ��c^���&Z�~t!��E��Sǌ����L�ǖʆ�$tܨ�t��� ^嶖��cx�>�m���f�t"��g}z�?(3�zM�6�;C��c:*g	�g�B �����z_��}2�����%�C�EMJ�$ȎO���i^{mM���E�-��5fέ�{gV��}+��.i�y�O�;����:�ćFm��M��ö:����aBy��~��Eu���q�-��!|�>�;�}|0�X| j ,���p�i�u�;�3�[�Q���z�F�\'��ತ<�f_6�h'�6������\����Aď���.��q�U �.����'��E�S~`���o>�9�|��|��!���(�2��-�i���J��KT\�U�	��K:��
��<�i&˝�U��u]�%��X<J����;E:I�O�����Cۥ]=km+k�c��F�u���������˜/�1]%�/��R��齌t ���/��%��0	͌a���൅,n5��Ѡ��5t��$K`/c,W�k����q�����B��m���ח��~G9�4��� �n7��Ѩ���;�~@���鿡�Y��i�6"苢���i�������֐��1��͌����U��CC#�t�6\�h�ؔcά�7���\g@
�����o�w�4������u$�tⷣ9�k��O�e(��Ɯ��``a�}Co������w�IA�ȲC���˪�M��g��Bƪ��d�U:����BŷH%:��t�f�ܔ:��'���$��P%!?;�a!&FUR�k-����u�-������'�Λ����4�Нt�v�|��i�k�o�� Od�8�u)�m�ɅuE����&4�����/�9Ο�[�sǚm�����E���,.>�#��w['�o�Z���Ybc��� �������@��U_&�C�u%��3��!R=�+�����n�w2���O��"��65��	��*��5���ש�j}ZM��Z�=a���jO���3'�Z�����5��`��� ��)D
��+�*�cT=�F_r��G9��)��[���c����;�P:o�n��G��K����B*t�ʈ��y�����8�����e�dt4�S���/T���;�	o+�e$�n�#{.t�Mc��x�h7�R7���y�k�̄��{�e��%�_'���n�f�9�"z������A!1�իY��ٔ��~:��29�!X��W����p���B!%�|�Md%3J���|��ʀ��D�ڍ�H��'�f�W�Z��s�����-����9a�&���5��b���B��n���[b����f�c�:������e2
�a6��}�D��945�?
%Ɵy�d^u�\`�X��[������d$]I��f�����{�[����)�x�ir32��59|�і��������޷����*�'8�)u�Х{X������$7rdM*��"���/ؐ�vLzsD����|#U�yuMB{K������ zx��}��[����Ԉ�сhY�E-i�(ٗ�ڠ�@۠I#l�iro����Ez����4���c�=�����c�]�]�lr�$���@���B?�w<z�����/�G����Ԉ�q8hno�J�A�3�l��9�"�A���g8��]4[������Ҕ�5ֿD^��O8�-��:nF�P���[��8�	#���9��Z5T�@]���w�W�T��.�|��eC�?)�<.qɠ$9��tl�u��P��A�t_�V��B��ĉsC�x�����b�B��ʸь2�*\��4�`���k2G:�ʱ�V�Ŧh����b�R�ˮ��g�30�w��Q��;ҒH��dv��	�a�A���3��Ɏ
��B�=�Gp�NF�?d¡P�G��Lƥ�'�ǌ�����<��
0�b�oV�E��WCC������
"��{�g����ς���Y_���*V����g��EEL%5(S|k���/0G��gw����؞����|�{x��F5�?cN�(��V�z�Ӈ�M�W���=�e�4���V��P1�N��7�7�V��/�_N�Zcf�a��a@��7l7�1�� 8�����E����q3ln���a@}7���>�Ei�o
|�8�����-s�'�`�`�]�U�����Wۊrk����1|:�q{�u�r�﫶���r�﫦�M�G&;-�QA���;��HZ<, ��	���B{�*�� �h�N�B��x{c�m�����Ճ4���>��R�(����ǐMn��S��q��n����ڊ�wK�}B��J�T�1�ۦ�E�ૌ��Z���K�`k���6�#t�a�ǒ�@\�ik+���Ngp�}���J% ��If���i���sV�̀n�+��u��3j��jg�[ݘXp<��Ds��/JO�Z��R=ͱ�Y]�q)\���H��p���㠽" ��1��~�i�
�l{
�A��xC�Ą�#G"�b�N��<�����!�гB���!,��U ���(ڗѼ֊
�	���bC1����I�&f&���毬5��"��Ҝ����u��c����rb˒9��lf��7�6N�;f�"C�ک���$Rc�}dl�{���\:�֓-�Ú������� ��*t'�BU5��.��ĥᖓ����LɎ�$�L�|DW�8�ZQ)s�.:��x� :n!�=��N	Y����X�T�Y$$����+���g�ϊ��қ�Zӥ�N���W�$�#�fQ�E����`��(������P<�����_<c�Ƥ@�������C3���Q�A���16kz
�i�Bh���&2 �YேBX0��賊�V���.��4_;#n�����"/��kJۆ�������L{\{s�+ރE��F� ���$���, ��ւY���E�Â��Yp�p�1hP3#�y�8����JF���%�S�e�~�yon�v��.ue�6mIb�1(cK���}|E���Fm0�_�3J6�21֎���VE�R�oa74�oR�41ց9Ζ.ɎoXdir̗�[�T0�_�'!�����H�5]iCc�'�_��O s��0h�y3VրԬ��i��1��<�2L6���h$伙�W��`��n�L��z��5�3@�����E�E����-|{~!�C�/i��b���Dƛ��׸�,/bd}B�زN]Ѣ�r��1�T�Ѣ���hs�8��b�O?�o���O�A��o���7����Yu���)�i�[�%�0�/1R�5�����Q�9�e�-��2c)g��\��6�����`�מN���M�]7{��|�\rߨ^����r������׾q�ڴ�߉	��j�<ʒ��m{ԡM�n����&���<��f��OQ*�E¯>�Y�Yc	��<�ó�4�{(\�!3�c�Xb�薷�񣅸�B��� "\�҆Q�������=�m��h��g�#4g�r�X��n����%�f���k��6TtQ3�E���>�Z����&ip]�/b!�a:1�i��I��~�i���J�"�����y��~�:sX�˄������`�'��~����M3�[s�Fm�b��8���	�����0�l9�q�FM':32��O���@o�~�����0�O�E,�f�,��i���mHT�6��A����c�@_����h�O��i?̓;3��ea!)R�E�Az<J]�j����oX�\�^���֔��\s1��.�@M�ю	�hR�mE~���]�~�
!�����U��r(ȶ���*�T���~��J<�Z�Z�S�M��!�l��\��V��ڀ��.�:c�{=�����9	�i��i7�F�\S�l�ST�~���n�8E��R��B;��-?����I;:m�"
�ܤ�j��������a�4Տ
�(^���:�;4�L�.k��Ly��C��\��k7m��/����&�,���:]����j�n{m�*��}���l��%���a�,x&+c���DfDF����gP��F��5B���km5k�ץM �t��+\�r�j����+�kF����Y�����2r����*��/��Hqu�H��E���o�� S����a�%��$ͲD3����SAx-����Q�Y1�W�G�*0��v�#s���s��<�7h���f��q~���H���\�������sRƂ��4a&u�S��{á�����c��s]�����S7�%%�u����j���c�����M������<�٤�Э�R���l�f�!e�f�j{�Z����ݽS���\#����n���]����Bb��Sx�!���� km�yB� ���u�I�~�m�b$�i2;�:뙫1��1g���b�	�g��e)���a"��S[���ݩ���z��)�"���B�`�٤�����c!�b�{������ޤ��jdS�b8����kz��\&�
����C�,�8��ޥ�O�&��`	�`�)���.�eKx�ϫwBӴ������,�ë�CͱwB�e�����&�Б��]��������������a>n�?��\�����i��O���0�P����Rѵ�����m�c�9&�Նe��jW|����C�Ŧ�b��g�p���8}��ǥ��X��圌N��h�kߤ`�e��`ź�ȓ�I����7���ڥ�#����Ó�'��D�dë�/kᶳ�� �D�U����$�l�@�����` �V������l��C`ŋ����R/�G|���� �7�ia��qb��m�ua��� �/ϩ���w|������l0#���o��n#$Ta�>�|m��������+�ū�,>' ��
�g���c��ݒ��;ή�]c�������$����ū��>'��5�ؠ�\ëޤ�}#$w;h6%���b�o�>x�w�>D���E�ݜ빔ޛ��e����H�d���(�y�M��\ƹ�a�H�3}��4�� ���1���ۋze���U���'�e<ζH�f��]|��*2�S���U���\��C��le�'^�� ��i\������A��$Y!�GsZ���7>�ZQ��^u7�I��A��3N2��I�M�
I9̮}�o)��Ǥ����̮����3;�4�q>�9i�s-;rd�$��ҁ{�a��hlY��ܓ��A��m_���Vǵ��$��K��[�S�/�s�"8��]t4�v�(0��~;�g"k�i���$��8��]4��!5@vmTV������삩��d��r��'lby/���Dw�Ť��sf�0��"��e��[ d��9(��sƜ��-b�1���]����?d��u�${ ��:�	&#o��b��(�����*='$�=g��f�}�̋��s�\*(��`�]�i�\*(�%�n�7�f����ą�ҡ������l���k��I��_��t��l�����1.��A��@��V��P���X�侚'�k�`��opa\VBS��C ���˅�勅�!%9�sëa��c��,�+���"��Ǌ���������k���
N�KR�Ьr��B
��h��('�y&C43ڦ�W������i��%�z[��2�a� <N�O��d��3M���j��7��l�.�b���$�NC��+����*��:n��k�L)�fe?�1�X5����,��HfR��0CÞ���M� e�Ah��NT2�aZ�جr���R�'�y�=' ��,�����b�4�a��$,�y�>',�'t��Z��e��� �,����AV��e��Ęk����(��m9!�@�:�$x�W�E}�Pe`�H�ka�ȑ��e�s,�����qCU�q0��`	�<�g�hX3���

��a��hS��d�E���ۇ��h���z�}f�$é X�|��nZ,b��Y!_$br��g瞃���W�W���ۜh�R��6�t�����;���0������U$��ǜ���55��X%`���gݵº�O�2��b�7��]�`�mX"���!ʨC ���
���a����<���=��'˯ ���|��ci����=��&�Ë���b�x���hݴhʼ��;�n�o!��ӟj�Z�����(�o? s;������)��a��������b�sO��?t6��7ʭ)�ML��J<,tJ