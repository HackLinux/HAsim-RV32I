;*�M*,-��-�;*�N*,-��� �Y��*,-��-�;*� �Y� �Y�]���_�_�_�^
���S*�S���~*�S*�O��*�S*,-��-�;*� �Y� �Y�]���_�_�_�^
���P*�P���~*�P*�L��*�P*,-��-�;*�O*,-��-�;*�L*,-���      7 �  $        +�WM*,���      E �  $        +�XM*,���      D �  $         �      � �  $  �    �+� �� �+� �M,�z� �N-� �,*�M� -*�H�[� �,*�N� -*�I�[� �,*�O� -*�J�[� �,*�L� -*�G�[� �*�M�z� �M*�N�z� �N*�O�z� �:*�L�z� �:,�Y8-�Y8�Y8�Y8	 �:
*�T��
�l� �:� *�T��
�� � �:�A� 8888	88	� >�?� 888	88	� �@� 8	88	88*	��Y:� A*�T���jW*�C*�D*�E*	�B*,�H*-�I*�J*�G� L*�H� *�I� *�J� 
*�I� �*�M*�H�{*�N*�I�{*�O*�J�{*�L*�G�{�      � �  $  �    � �:::*�T�� ��l� �:		� 	� �� *�T�� ��� � �:		� 	� �� 	� �:

�u:� � �Yc8�r:	� V� �Y*�T���k:

	�� W*�T��*�T��
�� :� �� � �� ��� � �� �2:� $� �Y*�F�s*�F�t*�F�m:*�F�s8
*�F�t8#8%8
#f$f8%ff8�� T�� M�� F�� ?*�F�p�� 0*�F�o�� !*�F�q�� *�F�n�� �� �Y#%*�F�m�      �   $  �    �*�T��� D*�M�w*�N�w*�O�w*�L�w*�Q�*�R�*�S�*�P�� �L*�T��+�l� �MN:*�T�� ��l� �:� � �� *�T�� ��� � �:� � �� � �:�u:� � �Yc8�r:� e� �Y*�T���k:�� W*�T��+*�T���� :� �� � �� ��� � �� �2N� � �� 	� �N-� #� �Y*�F�s*�F�t*�F�mNc8�s8c8�t88�� 	8	� 
n8	�� 	8
� 
n8
,� ,� �Y	
	jf
jfc8�mM*�T��,�jW,*�F�p8,*�F�q8,*�F�o8,*�F�n8-*�F�p8-*�F�q8-*�F�o8-*�F�n86*�F�s8*�F�t8*�C�� �6*�C*�Db�� �� 8fn8� $*�C�� 
*�C� 8f*�Df8*�E*�Bb�� �� 8fn8� $*�E�� 
*�E� 8f*�Bf8�� 
68�� 
68�� 
68�� 
68bb�� 
�� 688bb�� 
�� 688� #� �Y*�F�mM*�T��,�jW*�C*�E**�F�sff�D**�F�tff�B*� �Y*�C�Z�H*� �Y*�D�Z�I*� �Y*�E�Z�J*� �Y*�B�Z�G �:*�T���l� �:� *�T���� � �:�A� .*�H:**�I�H*�I*�J:**�G�J*�G� ^�?� **�H:**�G�H**�I�G**�J�I*�J� /�@� '*�H:**�J�H**�I�J**�G�I*�G*�M*�H�{*�N*�I�{*�O*�J�{*�L*�G�{�      (     � ��  � ��	PK
     �K;O�;#  #  (   sun/print/ServiceDialog$MediaPanel.class����   1   ! I J ()I ()Ljava/lang/String; ()V (C)V (I)V (Ljava/lang/Object;)Z &(Ljava/lang/String;)Ljava/lang/String; (Z)V <init> Code D I InnerClasses Ljava/lang/String; '[Ljavax/print/attribute/standard/Media; 
access$100 access$1200 access$1500 access$1600 
access$300 
access$400 
access$700 
access$800 add addItem addItemListener addMediaListener auto-select border.media cbSize cbSource clear createTitledBorder fill get getDefaultAttributeValue getItemCount getMedia getMediaName getMsg getSelectedIndex 	getSource getStateChange 	getString getSupportedAttributeValues 	gridwidth indexOf insets isAttributeCategorySupported isAttributeValueSupported itemStateChanged java/awt/GridBagConstraints java/awt/GridBagLayout java/awt/event/ItemEvent java/awt/event/ItemListener java/lang/String "java/util/MissingResourceException java/util/ResourceBundle java/util/Vector javax/print/PrintService 2javax/print/attribute/HashPrintRequestAttributeSet $javax/print/attribute/standard/Media ,javax/print/attribute/standard/MediaSizeName (javax/print/attribute/standard/MediaTray javax/swing/BorderFactory javax/swing/JComboBox javax/swing/JLabel javax/swing/JPanel 
label.size label.source lblSize 	lblSource 
pnlMargins remove removeAllItems removeItemListener replace 	setBorder setDisplayedMnemonic 
setEnabled setLabelFor 	setLayout setSelectedIndex size sizes sources strTitle sun/print/ServiceDialog $sun/print/ServiceDialog$MarginsPanel "sun/print/ServiceDialog$MediaPanel sun/print/SunAlternateMedia this$0 toString 
updateInfo weightx weighty  8 9 : ; < = > ? @ A B C D E F G H \ ] ^ _ Ljava/awt/Insets; Ljava/util/Vector; Ljavax/swing/JComboBox; Ljavax/swing/JLabel; Lsun/print/ServiceDialog; &Lsun/print/ServiceDialog$MarginsPanel; (Ljava/awt/Component;)V ()Ljava/awt/Insets; (Ljava/awt/LayoutManager;)V (Ljava/awt/event/ItemEvent;)V  (Ljava/awt/event/ItemListener;)V (Ljava/lang/Class;)Z ()Ljava/lang/Object; (I)Ljava/lang/Object; (Ljava/lang/Object;)I (Ljava/lang/Object;)V (CC)Ljava/lang/String; (Ljava/lang/String;)C (Ljava/lang/String;I)V ()Ljava/util/ResourceBundle; $(Ljavax/print/attribute/Attribute;)Z (()Ljavax/print/attribute/standard/Media; )(Ljavax/print/attribute/standard/Media;)V (Ljavax/swing/border/Border;)V (Lsun/print/ServiceDialog;)V (Lsun/print/ServiceDialog;)Z )(Lsun/print/ServiceDialog$MarginsPanel;)V %(Ljava/lang/Class;)Ljava/lang/Object; 2(Lsun/print/ServiceDialog;)Ljavax/print/DocFlavor; 5(Lsun/print/ServiceDialog;)Ljavax/print/PrintService; 4(Ljava/lang/Class;)Ljavax/print/attribute/Attribute; O(Lsun/print/ServiceDialog;)Ljavax/print/attribute/HashPrintRequestAttributeSet; 5(Ljava/lang/String;)Ljavax/swing/border/TitledBorder; _(Ljavax/print/attribute/Attribute;Ljavax/print/DocFlavor;Ljavax/print/attribute/AttributeSet;)Z `(Ljava/awt/Component;Ljava/awt/Container;Ljava/awt/GridBagLayout;Ljava/awt/GridBagConstraints;)V `(Ljava/lang/Class;Ljavax/print/DocFlavor;Ljavax/print/attribute/AttributeSet;)Ljava/lang/Object; c  d  &  2  4 { [  Y | Z | " } # } K ~ L ~ `  M � )  -  /  X    $  O  b  S  W 	 T  U �  � V �  � P � 5 � N � . � ' � 3 �  �  
 a  Q �  �  �  �  � * �  � R �  � ( � +  ,  0   �  � ' �  � % � 6 �  � 1 �	 f �	 f �	 f �	 f �	 f �	 y �	 y �	 y �	 y �	 y �	 y �	 y �	 y �	 y �
 f �
 g �
 h �
 h �
 j �
 l �
 m �
 m �
 m �
 m �
 m �
 m �
 o �
 o �
 o �
 p �
 s �
 t �
 t �
 t �
 t �
 t �
 t �
 t �
 t �
 t �
 u �
 u �
 u �
 u �
 v �
 w �
 w �
 w �
 w �
 w �
 w �
 w �
 w �
 w �
 x �
 y �
 y �
 y �
 z �
 z � n � n � n � n � MarginsPanel 
MediaPanel   y v  i 	  [     K ~    L ~    " }    # }    Y |    Z |    M �   `       �        *+� �*�*�� �*� mY� � �*� mY� � �*� � gY� �M� fY� �N*,�**� ߸ ��*� tY� �� �*� tY� �� �-� �-�� �-� �-� �*� uY��� �*� ���*� �*� �*� �*,-�-� �-� �*� �*,-�-� �-� �*� uY��� �*� ���*� �*� �*� �*,-�-� �*� �*,-��      +      1     + -� �M,#n� �M�	,� �M+�      k    7 �    *    +� �M+� ��,*� � v*� � �>� g*� � � \*� � �� ;*� � �� 0*� � �d6*� �� �� r:*� �� zY�� �W*� �*� �� �� q� �W� �,*