�x��^C�����x䙵�^���<^߆Ԇ��^<����<���������Fx���@A���-�������C<<<^^�F^<������@^�L���FF�F�F�F���������@F���A�AF���F�F���@��xF^@x�Z����fiyiiieiiyii��iiiiiyyyhyhhhyyyi�����������ūǭ|���������������pQp}�b`�{{�{{|��������[�rl�ll}b��}a}��zklzznaaQKZ������������������Ǣ��Œ�������j�f�Nfieiyyyiyieii��iiyi�f����]�yii��y��������������������������yyy�iii�N�W�������������j����N�e�eeiiydSydi�����������C����Ԇ�C��L��^^^xxF��x�x�x������E����������E��E����L�������LЩLF��x�^^xx^F�x����B����xxL�������^߆��<������<�����������<<���������x--�-�!@�;<<��^;FF��Ԇ����;F^F�����F��<Ԇ���F^���FF���@��F;��^���^��@FFF�^^Faib���yyyiiiiyyiiei�iiiyiyShyyhyyhyy��������Jt�ū�{�����������������Qa[[���{����|���||�{�purrp�����`�b��r}}zzzaaZ]]����������������������ʵ�����������f�iiiyhhiiiiii�eiiyyyi�����]�i�y�yy�y������������bN���������yy�yyyii��ff�W�W���������������ieiiey�lSddhi�J��Й�L��C���C��CԆ�C������x���x�������������������E���D�DD����������E��ʵ���x�x�^x�x�����B�ȆB^��L��^�C���߆Ԇ�^�<�����t�����<�����:��������F�^^F����^�^���xA�AF�F����B������@F^�F��xA�F��@�@�x�Fx^��Fn��N�iiyyii�yyyhyieiiyyi�yk�hyhhyyyl��j��������ūǭ�����������������[]p���|{�������{�����U���b�����|�����b[}zzaa]Ka��������������������R��ű�����{���e�iyihkhiiyyyi�iiyyhyi�N�`�K�yy�i��y�iyy��i����ibi�����������yhhhhShyyiff����������������f��ii�d�h�hghhi�J� ���^�C����BCvӚ�Æ^F�ELxx���x��䙙������E���������D�����D�t�E�𙵙�E�ʵE�x�L��xFxxx��^�ӆ^���^���J��x^���^��Ԇ����x�������������<���������<!!�!!!!�!�<������FF��^���^���F���xx��F�����;<FF@@^F���^^xx���FF��FF��x����AF���a���iiihyyiiihyyiiiiyyyyylSkll�llhl������������J�R�������������������aP����|{��Ǣ������������{{�|�|��|�|b��llzaZ]]b�������������������ǫ��㮝��������iiylll�kSyyyyyiieiylyHii����K��yi�y��ii�i�l���������i�y�yi�h�y�lzanznaz}�����|||{{�{{�{||����}lSSzzkkzkhy�J� ��xB��CC����C��C��^�����F^�x��䙵�������L�tD������Lxx�L��E��t�ttt������E����Lxxx�xx�L���xF��Ԇ�^L����^����^�B�߆���^<����������<<F�������2  5��!�����F����<�Ԇ<�^@�;^Fx���xFF�ԆF@���<AA5�F��^�^xx��F�^����F���A�Fx�xA�<z�y����yly�iiylhiiyiiyhhllShkzklz�ny�����������ի�{|�����������������bQ[���|��{{���Ƣ���������{||��{�����b��}za]Kp�������������������������Ţ�������yll}lzzlgllhlyyiiiiyyhyii���[K�yi����}�iy�i���[����}�����y�y�y�ylq�qqqqUpp[��b������������b�[UaZZZQ]Z~]ZSij�D �������������C����^��x�x���x���E���䙙��D����t�t���DD��E����D���������������x��x�F��^x����x����x�^��<߆Ԇ߆����F������������<���������F���:��<<��<<<^��<����x��A��^��^�Ԇ��FF�����L��F^�����A������^^��Ԇ�x�Lx�^��xAxx�����xn�y�yyyyhyyi�yhyyiyiiylyhlhglk�kk�n���������t��J��{�������������������}Ubb��|��||��|�������������������������zq]Q�������������������|�ǩ���ܫ�������y�kkkgkhShlhyhiiyyiyh�iy�i��p]l�i���}��������������l������y�����lzaaaaU[��b��|�{���{{||||`�b�}zanknn�aznSyW�D�tA�B���C�Ȇ�����C��^�x�^x�xx�E��L������D������t��������^�E �����E��t�E��������L�L��x��^߆���^Lx�^����^߆��ԆԆ^<�^x�E���������<<�F<�����������^^�������������F�F���^�����@����^��������FAF^x���x��Ԇ5:x<<��A��F���F��F�xx�A�^�����A�x����x�kyiiiyiyyyyyyyyyyy���yhyllhhSlhlkn�������ǫ���ܫ��{��������������������}[��`|����`��`������`�������b�����b��}aQY�|�����������������������Ţ�ʫ��{����n�khhlghllhh�y��yyyyyyyyii�pK�i������������������i�����iyy�i��yyhhhhyyi��������������������fiyhdhhhdyhhhy`�tD�xB��B��CC��Ȇ�B��߷x�����䙵�����E�����DD���v��������vvv���  ����������������xxLLx�^^^^^�x��^�����^^�Ԇ���^����A��������<����������������:��<<<�<�<������������F�xx��������^^�FF^��Fx�xxx�߆��AA5F��F�@��@F�����F��xF�F����A�xFx�kyyiiiH�yyiyiyyyyiiyyyyhyhgh�hglk�n����۫�����D�ʫ�{�ь�}���������[[}[��p���������������������������������[�}ssu�pp[���������p}�����ǩ���Ǣǩ��Ǘ��l��klSlSghyyyyyyyiyyyyiyiii�rY���������`�����`������������������yy�yyhyi�f���������������j���HyyHyiyy�hhhh��tEx^�ȷtL�BC�C�^^^�^^x�^F���������E������뵥��������������������������?tt�����ELx����L������BB�C̚�^^xxxF��F^^x�A��L�����<����x���x����������F�^�^������F�����x��xF��^�Ԇ�^^^F�FF���Lx�@߆�@�䙙����FFF�F�<�����A��F�F��x������xF�x��kii�i��i�yyieiyyyiiyiyyy�igShShlk���n��{������ǒ����}�}������_mXooIo�cw�r����}}���������������}}}}}l[}}}kzzZK�ww�~oo~oX�_�m�������}�|{����|�����]knnkklghhhleyyyiyiiyyyyei�ii�r]��������j��{����j�j��j���`�``�������yy�yiiN�f����������j��`W�NylzSiieNieil�lN{Jෆ����LxR��C�����x�xL���xx�����E�������L�������W�W�WffW�f�����bu�� �L���tE��������x�xF��F�xx�B�C���������x��^^��FFFx����x���<����x�����������E������F�����FF����x�����������:��FF^<�B��FFF����xx��xF��^������xLxF�����^���x�������A���F�x�Fzyeiiiiiei�iy���yyiieiyyyyyhhglSk�kk�c٠�i�iiiii�lznmO�k��ߍ__g�m~~YY]cw�qzz}zakzl�l�llUz}klaaZnnazazzzZznn~��wwsmYYomn�g_m���gOmnzzlhii�i��bǅszkk�khhhhhyyyyye�iiyy�ey�iii�pQ�������������{������{�{��������`���ii�i�N������j����{�j````�N�lPsQiffWfNNlll�|�x��B��BB�xLx����FxF���������������D�L�ܥ�r����W���aqq�uqr}N�fW����u�J�Й�t����������x����^^Fߚ�C�����������^����^���@xF���F�F���x��������t���߆����^��F�xx���������������A��F߆�BB������F�x��F�B�^��:�x�xxF�F^�^�<�^F�x�����������FF��Fzi���iieieiiiieiyii�y��yy�yyhhhlkkkz��yyi�iiy���lnn�gn���m��gnooYYXcw�sqZannnazzzannnnnnZZZZZnZnZn~��wwVoYYomgg_�m�ô]kkOnnkzzkkkllhylƹ�zkkk�lhhhyyyy��iyiii�ieiii�f�rZ�`j������������{��������������{�������[��[�����N�`����bbbb��[zUQs��W����N�}}�|�������B����Lt�xÆ�x����൙��E���D���ʏu���fWW�aqq���������qr[N���������L���E��൙�L�x��xx�x���C��BB�^�����xF�F���^��FF�<����������������������������DDL���������������������t��������F�<����^F^F�;�xx�L�xF�B�x^<���FxL�^�^;F^���^��x���^�xA��xx���xFPle�fiiii�iiyii�iiiiiei�i�yyyyh�kkkk~��}iiN�jj�`����nnn���mm_���Y~omTcwws]~nYm~mnZZ~ZZn~YYZmZ~mZ~~n~~Z~m~��wwVXo�~m��mmm�ߴ�nnnmn�l�iyy�iiyl|�c�kkkklhyyyi�i�eiiiiii�iei�f��rZ������������{���{���������������j��}zanaaaUaaUUU}ppppUUaaPPaPZnQ�Qb������b�������ӺC��߆Ԛ��LE���x�x�������E��Dtx��u[��f��[uq����������׶�}q��f�������F����������xxx�^���ӚBxB�������xx��F������^���Ԛ���������������������������������������������������    ���^��<�^��F�;��FxxF�^����^�F�xxF���F���;FF^A��<�Fx���x�x^��FZ}iiiiiiiiiyyyiiiy��ieiiyi�iyhhkkggko��li�������j�j�zn~���mmmmmmno�YYww�s�]YYYm~~~~~YY~YZ~YZZm~kY]~Z~m~~~~�\�wwsX�oYmmmmmXrߗ�nmmky����N����i`�ckkgkklhyy�iiyii�e�iyii�Nf����qZ�����������{{��{{{{{{{{{������{���}zZZYYYYYYYZZZZPPaPZqQQ]Q]]QPQs��`||��`�����B�C������^���F���������E�x�E����L�ܼr��W��������������������׽�}\pfNW����D���򵙙���xx�^�xF�B�^Lx^^����������<��������Ẻ������Ӻ�̺�������������������������������������������    ����;�����^��F�F����F�^��F���x�������F<�����F���������Fx^<F�FQziiyyyliiiHyhyiyiiii�iieiyyyl�kzkkSV��yi����j�j�����nn~�߹XmmmmmO~~~o�wws�\Y~~m~mmm~Z~Ymm~m~~Z~nY]~Zm~~Zm~Z~��wwsX~~mOmmmmm���nnnz��`�����������sgSkkkz�hyyy�eieNiiiyiie�f����PQ}���jj���jj|�bb��������`�`�`��b�[pPZQY]Y]]]]]]QZPaUaaPZZY]]]]YqQ����Ǳ�ј���������vӺ����^��߷�E����������E���p��������������������������ױ�zZ�����������xx�^��^���^�xxx^^^���x�L�x��^�߆������ӹC��ȥ��ϏϤ������޹��ں�̺��������̺����������������  ����^<^F�^�F�@��FxF^�^�����x��x��FF�FÆ��F^FA������<�F��^���F]ayyly�yyiiyh�yiyhyliii�yyhhh}��zkkkc�jyi������j�����}no�߹Xmmmmmm~Ymocwcs\K]]~~YZZZm~mZ~YZZ~mZYYY]~~Z~Y~YZZ~��wwsmYY~mmmmm_��ȁmnz�����jj���������lkz���lhhhyiiiillyyyiy�����jP]}[�`��{{{|`b�[�[���b�bbb��������}aZYYY]]]]K]]QZUp[[[[pUaZQY]]]Qq������ũ�������Ȇ����C��̚�Ԇ^�F�������������낏���jpa�����������������������Ľ�Zzi���ut�������x�����^^^^��߷�x��x�L�թ��x���߆��������ј��٥���ҥȥ�������������Ϲ������ں�����������x�  ������<��^F��@�F��F�x��^��^F�����x�x^�^�F^�<FF���A���A�A�^^^F����F�]alyyyyiy�y�hyyyy�iiiyillhhl}zp�zkkzcٌyi�W