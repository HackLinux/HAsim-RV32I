 T       l      U       T    T   l   T   U    T       /      �� ��D����  a�  �D ��� �������         M          ^   �       ��� p�D����    �m� p�D ���=           �  �       r  �   q   
   q               M        ^        �    M        M   ^    M   �   3   �^        ^   M    ^   �    �        �   M    �   ^    2      �C ��D ��� �D  �D�������� ���         �          ?         D p�D ���    �D p�D����r  �   q   
   q           ]    =           �   Y   �    ?    �        �   ?    ?        ?   �   Y   �:      �C  aC ��� @D  �C���� �������      s      �     t         �   	q  �  r     q         �  =      �      p  �   o      p    y  )           �         q   
             s         �  !   �9   �   �e   �    t   W   �   �       W   �   �    �  W   �s         s    �  !   �9   �   �e   �s    t   W   U   �s          �s    �  W   ��      *   ̧  s     �  t    �     W   f�  �   t          A   �t   s       U*   U   �t   �  !   �9   �   �e   �t       t   �     �*   �          U*   �   �   s       A*   �   �   �  !   �9   �   �e   �   t       �  *   ��       �  s       ��  �  !   �9   �   �e   ��  t      ��      =      ��  �C����  z� ��C �����������   �                          ]   v  �     q  p  �   o      [    	   [              �           U   U3   U=   U�        �            �    %   U=   UL   �   �   �               %   B=   BL   �   �   �   �    *   �       *   �      %   L=   L   �   �L   �   �    *   �          B   B=   B   �3   �         L   L=   L   �3   �>      HC �mD ��� ��C  �D �����������                 �      �       �TC  }D����q  r   �      ]    =    
   q                              �        �           J   �f   �         �       �          J   �f   �        �      �    �       J   �f   �       �      �   �    �        �       �      �   �    ?     ��C ��D����  �C ��D���� ��� ���         2          a       ��C P�D ���q  r   �      
    :       v  ]      
      
  �            2        a    2        2   a    a        a   2    @     �"D  z� ��� @5D  /� ��� ��� ���   "                S  p    �  s   q     q      [            	   [   q   
         "       =   U
   �   �"    S     �9   �"    p   =   f   �   "       U   U3   U   S     W   p      �9   �S  "       �S     
   �S  p      �p   "     p       p   S   F     ��� �(� ���  H�  � �����������       n            �       @�� �%� ���    �T� �%�����   [   )   p  o  �  p            y  p      n       n   �       n       �   J   ��   n    �       G      �� @� ���  HB  �� �����������   �   d     �      	              B   �����   [   )   p  o  �     p   :      �    d    �    �    �    	    �        d   �     d   �    d   	    d       �   �     �   d    �   	    �       	   �     	   d    	   �    	          �        d       �       	    K     @5�  �C��w� �(� ��C�.����w��.��   Y         �      �              ]   �     q     :   
      [    	      s   p    [           p  �   o   :   �        Y        Y    �   ^   �Y    �       Y       O   �   �   �      �   �    �   Y       l^   l   ��      #   ��   �    �   Y       O   �   ��         l#   ��   �      �L     @5�  C�n�� �(�  aC�]d��n���]d�   �     �         �        v           :   
          [    �     p      s   p       ]   v  q  �  r  :   �        �   �      ��         f   �G   ��   �      O   ��   �    �         �G   ��   �      Y   �   W   �   �      �   �   %   KJ   KL   Kf   K   �M   ��   �   W   ��   �    �       M      a� ��D ���  /� ��D���� �������         _          /       �;� P�D����   ]    =    q  r   �         q           _        /    _        _   /    /        /   _    R     ��� �	����� ��� ��� ������� ���   ^                 {       @�� `�����o  	   p     )   �     ]   v     p   :      ^       ^       ^   {       ^              {   L   �   ^              {    {   ^    {      %   {{       T      �C �"� ���  �C ������ �������       *            o        @�C `� ���p  o  �     	   [      p   :      
  
   
  �        *       *   o       *       o    o   *    o       U     �	D �"� ���  D ������ �������   l     �            *   !    �D `� ���o  	   p     p   s   :      �     [   )      l   �    l       l   *    �   l    �       �   *       l       �       *    *   l    *   �    *       V      �A ��C����  �B ��C������������   �     q     �       "     B @�C����    �  v     �  =         �  Z      �  o  p   	       )    [    :   �           q       �   q   �   �    q  �   d   �   �q  �    �   �   #   {   ��   q  #   �Y     @5�  zC��_� �(�  �C��w���_���w�   �      �     K              ]   q  �  r     :   
          [    p  �   o      s   p    :   �        �    �   �    K    �  �     �  K    K   �     K   �   Z     @5�  �B���� �"�  �B ��� �������             �      #     2�  �B����      ]   q  �  r     :   
   ]                [    �     p   :   �            �   �        r[     ���  a� ���  ��  /� ��� �������                        �     q     ]   v     y  p   "      @              %   fL   f          �e   �        L   f       L   �   �          {Y   {       %   Z\     @� ��C���� ��� ��C������������                   �   $      � @�C����    ]   v  �     q         [    p  �   o                  �               �    �          �   �L   ��         {   �%   �J   �L   �f   �]      �� �(D����  �� @5D ������� ���                     s   v        �     :      [    	      v     [                        �3   �          9   �U   �    s     �9   �          �M   �         rM   r9   �U   �   s     rM   r   �9   �                      �   s     �   �s       s        �3   �s      ^      �� ��D����  �� ��D������������         /      �      �   %    ��� 0�D����r  �   q      =    �     [    	   
   q        [                  /        �        �   =   �/        /   �    /   �      {=   ��        �   /    �   �   =   ��        �   /    �   �    _      /� ��D ���  �� ��D ��� ��� ���         �          M   &    �	� 0�D ���   ]    =    q  r   �         q           �        M    �        �   M    M        M   �    `      ��  zD ���  �A @�D ��� ��� ���   v     �      �         '     HA ��D ���   ]    =    q  r   �   
   q           v   �    v   �    v       �   v    �   �    �       �   v    �   �    �          v       �       �    a     ��C ��D���� ��C ��D������������         ?            (    ��C 0�D����q  r   �      
    :       v  ]      
      
  �            ?           ?        ?               ?    b     �"D �sD����  /D  �D������������   x          �         )    �+D  }D����r  �   q   �  :   p      p    y  ]              v  ]       x      x   �    x         x   !   �e   �  �   e   x!   �     !   {e   {�   x    �     e   x�          x   e   �     e   {   �    i     @gD  �B ��� �sD  �B ��� �������                    *    �pD  �B ���q   
      q  �  r  =         
      q         p    �  :   p      �  )    �                     �       j     @5D  �A ��� �AD  �B���� ��� ���       P              +    �>D  B ��� q  �  r  q   
      �  s         p    y  
      q      P        �!   �e   �P        {e   {   �!   �Y   �   P  /   �          P          k     @D �	� ��� �(D  ������ ��� ���   R     Q     "         ,    �%D `� ���   p   s   o  	   p  :      �     q         [   )   q   
         R   Q     �R   "    R       Q  R    Q  "    Q      "   R    "   Q     �"          R       Q     �   "    l      /C ��C����  aC ��C������������   �     X     W     q  -    �TC @�C���� �  r     :   �     	   o   y     s   p       �  =   �   \        v  ]       �        �   X  ^   ��   W   �   q   X  �      �M   �X  W   X  q     {M   {W  �   *   {   �W  X  ^   �W  q  *   �q  �    q  X  ^   �q  W   n      H� �"� ���  �  � ��� ��� ���       _           F   .    �"� `� ���   [   )   p  o  �     y  p      _      _  F       _      F    F   _   F       o     ��C @� ���  �C ���������� ���       T            k  /    ��C  � ���p  o  �     	   [      p   :      T       T   k      T       k   k  T    k      p      D  a����� �"D  /� ������� ���      S     @              �  s   q     q         	   [   q   
             S        @      �          {
   �S        S   @    S         {
   �@        @   S    @                 {   {3   {=   {   �   S      {   {   {3   {=   {   @      �   �3   �=   �   �q      D �(D ��� �"D @5D ��� ��� ���   
      w                   v  �  :         p    y     
    w     �%   �L   �
       %   �J   �L   �f   �w  
     w         
    	      w  	   �s      �C  C���� @D  aC���� ��� ���             :      �  0      D �"C����	q  �  r  =            q      �  s   p      p    y     �  )              �         q   
            :       �   :      G   �:   �  G   ��      �  :    t      �C  �C���� @D  �C ��� �������   :                 1      D ��C����	   q         �  =      �      p  �   o      p    y  )           �         q   
      �  :   q     :       #   �   :     u      HB  �B����  �B  /C ��� �������       p     �     �   2     zB �	C����   �  v     =   ]   o  p   	       �  )    	   o      �  u   s      y  p         q       p  �  G   �p  �    �  p   �  �    �   p   �   �  G   �{      �� @����� ��� ��� ��� �������       R             3    ���   �����o  	   p  �     q     ]   v     p         R          R    }      ��  �A ��� ���  �B �����������                   �   4    ���  B ���       ]   q  �  r  �     :      [    	   ]         [                        �              �    �         �   �   �3   �=   ��         �   �=   �~     ���  zD ���  �� @�D�������� ���   t               �   5    @�� ��D ���r  �   q   �     p      [    	   q       
    [                 q       t       t   �       t       �    �   t    �      =   �      HB �mD����  �B  zD ��� �������         �          v  6     zB �vD ���q  r   �      ]    =    
   q               �        v   �        �   v   v      U   �v  �    �      /C �mD����  HC  zD ��� �������         >          �   7    �;C �vD����q  r   �      ]    =    
   q               >        �    >       J   �f   �>   �    �        �   >    �      zC  �D���� ��C `�D ��� �������   >                  8    @�C ЄD����q  r   �      v  ]    
   q           >        >          >             >           �     �D ��D����  D ��D ��� �������                  2   9    �D 0�D ���r  �   q   
   q           ]    =                  2             2   Y   �2        2      �     �"D  �D���� �(D `�D ��� �������   b                 :    �%D ЄD ���r  �   q   �  :   p      p    y     ]    =       b           b     �     @5D  �C���� �;D  �C ��� �������                  
   ;    `8D ��C ���    q      �  :      p  �   o      p    y  q   
                    
             �9   �U   �  
      �9   �U   �
        
      �     �mD  C让� �sD  aC��b�让���b�             "         	   q      =               p    �  :   p      �  )              �         q   
      q  �  r         "     O
   �       
   �   �   �   �   �9   �U   �W   �"      G   �"        �   �   �   �9   �U   �       	   �G   �   "     N	   NS   N�      /C �(D����  HC @5D ��� ��� ���                 r  �  <    �;C �+D ���q  r   �      v  ]    s               q          r      �   r      r  �  U   ��      �  r   �      ��  �C���� ���  �C������������             =             ]   v  �     q     :   
   p  �   o      [    	      s   p    [           :   �           =             �=         �=         �         �   �   �3   �=   �   =   *   �      �� �"� ��� ���  ��������� ���       F             =    ��� `� ���o  	   p     )   �     p   :      ]   v     F          F    �      HB  a�����  �B  /� ��� �������   	      o         	   >     zB �;�����p  o  �     	   [      y  p   @   S     S     @      	    o   	    	    o  	     o  	    	   	     	   o   �      �� �� ���     @��������� ���       d     G         ?     H� ������   [   )   p  o  �     y  p      d  G    d      G   d   G          d      G    �      HB  �� ���  �B  ���������� ���       e     	      G   @     zB �������p  o  �     [   )      p   :      e  	    e  G    	   e   	   G    G   e   G   	    �      /C  �B����  HC  /C���� ��� ���       g     �     p  A    �;C  �B ����  r     �  �   :   	   o   y     �        �  )       	   [      g  �   g  p   �  g   �  p   p  g     �M   �p  �  W   ��      /C  a� ���  HC  /��������� ���   	              o  B    �;C �;�����p  o  �     	   [      y  p   "      @      	    o   o  	     �      zC �	� ��� ��C  ���������� ���             y     j  C    @�C `� ��� p  o  �     	   [      p   :         y      j   y      y  j   j      j  y   �      D @����� @D ��������������                 U   D     D  �����o  	   p     p   s   :      �     [   )      q      q   
            U    U       �      �A  C����  HB  /C���� ��� ���       u      �      E     B �"C����    �  v     =   ]   