�5������AD��a��,��쁛!�Ě��=�hxڎ�a�}q2��,�ZA�ɽ*���'�^��D��������
&[�Y�]Ht��d�u�;���v@f���}��*���*�"1�n��5�T Ms0]�2]���:��:s`�/�A~�cu�62�fR� K��B;Cw�Č4Ewz~z�ߞ�(������:�9M�1����/���9�)Y����:J�O��o�>�I	�rM
f2��_���c���.����_�%?�(�ҙ5���,��B�O�
<�9Zہyq0��c7�Y�	��z�!�:���܌
��p;���gP�ÎQ�$�N�ɋG���z4T}�I���,��ׯO�6�]���q��Jw(Q�|�*�کȴ8-wR�z}}�[��	D~���[�R;(yi�w�;S@:��:/��4y��X՗���}3D����R|�K��	�x|tؚ�?�S���&"MV�{SN��1��a=���}UI�9m�ol�T��z��-�C��8��4ŧ�Pڇ�|KU˭�J�\����~Wx�"P��$w�^�gQ��E�<9��n��2�ۂ�j���9 k�!T��r�
��E�⨱��>��A���ru���������5>��3o8������r~f�8M��3����#�a�l���d
����m����,D���+f�8���$.I�Đ}�T�}�3�ӡ�Ɉ�E�8Õ^8CLY��C�04NtK�V@�
�e�R|
1
�pM����]�_�h*й}�*�q�ZᏞP�{,�OF��>�V�^��}mJ�?�}�x��W;$x�M���&.C�7�;�z��2��=_�'���5�p~fm9�q������}|.34Uzp5�}0���}�>��3ë	�k�6Ig��6�}������ݠH�8w&	�Q��FM��q7������큜x�1"5����k�bs�^Wc�� �����_�'�!l���X� 4e�u���Mg&�ҽ� ;�^B���p���s����U��h��d��Q���d��tv�o��+�8|�УU��t&q�j��T�,PGT�M���5m��O��%	�Y��jl�t6��@�{+,pF&�z�8-!'[��-�'$?�-�Y�<p6��H�֋����{5��]0�7�v�}�H�"�lL@���*J����C���~�T�o����V;$4�$��jj������V}�K��7p2@[����{�M���*W���F�}%*�l���6&U�j/���j��{�5B��{��s;J�^l�0M���<�Ī"=�����h�c���!�� �M�s����kg��6�:4���]64e�
v*S˷5�I �Yc
_�'	��~��C�s~��bv��!��t��*Q�p�$1��I@�/���k�D�v��������ѓZ��� ]�/�}��^�����d�S��-���;�v75Bzox���e1�0A��{n�qS��I=��KʒL�oN�����~8C>�VW���kgC����J���Q�S���rf��z��Y��Q?�=���$��E�Kpb��/`�kK�	����{AH͎i�U\�����f�S�W�Dr5��{�S�8�1��Vd[[�a�!#=��;�N��y,�P�gXrf��!��>��� ~'���"Q��_%w:`b<᭤���]�