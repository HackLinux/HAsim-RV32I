-9999)_� Ns_I\~�#,PNA\���A<_�I��#, Az�8�� ,�1�,,5 5)sߌF&�  I<&N&1=-F���8�#�_#%,)N#,_,, s,\PA8" 5, I_AA8!
PAA<,,,5AI 
 5I<% \�sF_)<r�Ij~�˧_,�]<<\_FFj�,,sN�r,��s˗����A#s�z?PƵ _?, ���ٌ�5s-FFF9=<#\�\\sٗ�#AsNA���,��5�٧<AI\ٗ�1"��!9-#r�A%%A�,#  <�=9-FF#�5
��8bs�P) A,,,sP8b AA!)!8�##P AA%,#!,
�rPz,__�P,I�85
,A�#�<,j-__\��,����_���r\NP�_ \r�r�z� ,)�r�5"b�
,_FNF,?&_#�%_~P�r\�Pr��,PNrͧI���,N I��I 11P58Arb,z1FF--)91~1=jz AA\��8%"P#Ir8
% "%%8%�%%#AA N,#%#)# %��<F),�NN<\I�/A��,A,PI �,%\A) ,��,#��__��rN<#\Ʊ\_�I,s������쌱��,
#NNz� ,N_ _�)<, �˱\N�_NN#
8ƌ�""s,\\#�߱�sNP]T/%), /8 �jF��1-��=--z\NP<P �����]A�%%%5I   /%%)5
]T�A)A AA�_�#AN<A55��NN_�,_Fs,�A��A�r�_s\P � ƌ\����?&#\��TPsbI8,NAs��I�b5b���P\��� 5�s,_Ps�r,As��#\�#IN1)N�)�ƌ��zA, ˗�jTs��8T%85\8)����_j# 1F--j11�P,,"�"�88�\_T5�sA, 8],5�5
)#PP�5\#N< _rr�<A,�s]_NA]�,_�z��������,Aj#N,I<�A��_ss,��5�
5 �\rss5PT��Ir ��_A I,�sArs�� N5r�PA��)jF�%\��5\sAN&AN<,_z-Nb�5\5P5",,IIs���NF~~%<-~v_�<j)]//8T�IA%],,,�/5
IA �TI,�
�)PN~<IA \N,\<_A_A�b�#\,\\�\_z�~�#������ٱ�_�,�
 5/8 ~\Nr�IP#),s,\rs\ "T ����\s��P�s�s�#�P\II�,\�P,<#_
��)I,, \5#)�1 8�TI%r_%5/5�%�1)#< ����v�N11)%88"I\<55A �\
8%%�%r�I,A% ~#I 5r##NA\s_I)),5�5rs, <I#5�A�INN~_r�I����])< Is,�<#PrA?,A,\A)sI 5s%A�8I8%%b�,r��AP�A) A_�s��%%IrA\���,  < \As)s<~9-_FA5� #85T5A<]s/
, r ��_
T8�_Nz)I#]I%srr,�\
I58,,"%I5I�  %A\]s\AP\8A%I,5IA5AN#��8%��<)s_\)��T5 < Ir]IA5,�_N5#�A#A?A_r,I5_,\rs\88
8%\s,A\��,,<AA�)_NI�%,\��r#<N ,I,A\F)v)1F_��#,N/%,5s/#PIA�_)F)FF)/��1NI)�8"5/55s5/AP�,,5 
s8T
8 58%b,,58\\A)5A<<%5)<,#)#,I\%�#\__���]]%�r�%%\�A,_�A#_\AP�r,, 5� \rA58A
5sT%�AA_]\IAr,rT%�\r A, ,<#PA~
  �9_Fs\j&N�]A�]\<)I 5
%s,#��� I~�,,A#s,<�vF\_#8�8"%%AI8T]"A�PPP�<88"%5//sT%/#P)%

/A,%%,\P,)<_<#�,�Ir<~�A]s#�,Assr%5s�AN��P5s���P, ,P�,�\sN N_%%I%As\�INII
!
\P,�8s\P,\_ \�Nr,�I


%s~zP P)Is��)AA#_ 5%\)��,,,,�~8�_˗,AAI,A,~\jI8%�]%5]/5,ss5%% "%I\5I8�8
"_,)
 )%
)\I, ,P#NFzz_I5
sI� /5A� _\,,�\"r%I5��s\r%\rr_�55N_P\ s/%I%�5rr5%I55
8I,<\P,,rN,\ #ss��PsP 
]5%,\�%�#)FI�)),5%A]5�T% �� ss��#8/z�1%A���A\bT%8/T"85%,PI]/ 
8�I#<)
%<%
A]%%,PAN)�z<<~I]As,AN#As _P Is5, �P<P ,5P��s\sr,N##N,!A8%�%�s��As\)
)%5r%#N,<\,��%,�]%!T]sN,�#\ As) APr�s�\�)_˱\8b�5)1�z)%
]\�)I~5\\Ab""]%/"%<\�5T " �/
,N)#A)]Ir,\,,zsA,rAA_r,,,AA_N_\]
,I#�_I~_,PN,I,A_%PPsI#  \%#\%T%\��]��s�AI%A)I�5
IAAAAs5 ,P8\�A#<
%I#  I<< #I�<N�r%�
s_I�A�58�<)Fz~]#)\_A]T��b�5
�"8T/
���5/!
)%//8�

% A#A)A %%5]/"5]~_~Ns,#INP) s\r�P  5rsA5IsI_rP,%A55A<##5,\5%5II�P,5r5,AIs58T55NAAs55I "r,55����)\ #v%\I<)N# )~v<-_1,N�I8sb
�\\,I5\b�j1)z�A),I%II\AII]�8s�8�s85s��I5
s5
%88
%#A

%ArrI%rI58A\�<,\ )<r���A,,)AAI%5,, <rs\5%5 ,  NIA#)#%5Ab8%58T%
#�\A
I#)  \�~PII])N##_]%% 55\,I#,�,_A#\,,�N�\A�&9)z1F)#A��!�I%�ArI8
��FvvI\,)I���I5sT\�5ƌ5�% �5Ir���,))]IT55%\rrT�I) I
II5)5%P\�r<�\ T�A��A,#N<#) 5\I% sNN,I\55A ,,, 5]IA<#Ib��]\5A<_I,)_N#ssr\<\�)<II%5I%P ,PPsAP%�#~I%P�%�~))N#
TI�T\8�I�r]I58I%I�v9F)###\)\�b�8!!!I/"b���5<%A%
II�\r5)9/b%,\�T5�5,)#5%%s_5IA_,,Ns�&/"�P�sr\A<,,,5)IA%,s�N  %I%])N# #PA#%II�]IT
%TII)#,5I~ I 
,~<#,#)#,,A%5P#5,\,A<A%�%!rs5)�,<_NA�A5�\ssI
Is���)9-�_ #IAAII%%85!AI]]T"b�5�5]5I
55\I))%

"T8),,�8)I,#%
5%%AA% #ANss\r\\A%5\,#<)5)A� ,,\)r%s<#<<%I5
8]85A!A\��%5A%!�s#]))!<AA%r\,),\AAIP_�A55IA5%s~zN<_�r55s\�))<~r�\��),�#, A,)Ib
5T��T]TT�r8T5
%%)##\)I%"!55
)A\5*E4.E^ww���^��ccoo�;c^EE0a�mMU�|ULB�m66omaU6oLLBDo|||6$''B[LUMM'6mB;MMm��Mo||La6^n0.^^c|oL'$L|�L7*CCS^�oQ}}SGG*$*7^Ec[07*$ElSS}}GS^S�wLGeS00E}n0.[|��hha�|QUBamJXXh��m�X6XX'D6$$.LcUUaMo|��o|[;.[|UM6'.UoQQELLE^w�**G00xo$6$^�EGC007E0S�^nL.$^^EwwGSwGS}w�w0GS0CGw��E..LMhUDaLD;.DaD6JahJMDMmmmD'DXJ66';7'76..Ma�oM..o[BM[6BLMB.Bc}[7.$ELUU��cE$$$707E�lE[^c}�EGG��wEw}70C*Cw7o���hm.'6XaJJ6h�{JDm��a6'6'M(;'.6''Um60$;���o|M.M|M[����[7$6UDMm�|[.LM.;;7E^Q;.Y;00E}}c}�xQG^S�wE^}n^G*CCC**0$;�����a6B'JXmo�mDm{`hD66aaM66'o|aMMDXXh6[��oB';7;[Moa;oMa�����|;Dom|�������M666'$.$;L;;70E���Sn^E^��w^}�nE}SGSGC000o���|��aam6D6'J6.6DDX66DJD'''''X�MDJJDUU;.XX.oo�|MU7L(BB6.BMUM[M|��||����oL�д||�m6$;c;MLc}E4E^SLBL;}�����؟GwqC