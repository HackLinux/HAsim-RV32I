��y�)�~��|���-��3�k����g��Bz6g���i��s�0�5^���G�g�ޢ�}�y�3����g���8��gg��	���>{חi\6���I��2UL%���k�9�<Q�������r�ˎSan��v's�3�Q��9_8��!���� �/�$틤sZ�6�����dE�0jw���ڛ�܍��5
$��\���$��<�g�:��q`Pץ2�a��c��#j�Oj�N��4����5!����Y�oSOڻX���5����K��c��kz��C����yΤ�Gɶ3�/
�	�u����x���T��6����[���|�g*a㺞'wZ����JCG��w�də�`ik��.Scע/�n��y.���ذT%P�1L1u`���D��8ѦːqO 	��6NfWh�-#|L��˽��&�߀�p�t�}�`�-z ��V#���N�#���y�K2R�}��C4�ޞV%;b���=$e�n�$Φ�BԳ	��k.�HG�'
���V݇x�sD�,�VU�=�'RwꅰZQ����q9��!�`8�y6����YhӇ���D�֤��������9XCDS-��K.�zCdZ������a��λ'�A�Sl���׌��������W�{K����Q�U~��������l�5���9����;�r��{�ɺeر����Μ�I�z�~wJD��N�cdu� ���"��ٖ+F"¹ѩk|�h�O�\oSK�ڦΥ�N�i7��5�k6��P<Y���Ӗ�]�ʥ3X�C#�s�3��ޖ�w�Z=Z�n�[h#���x����]��T�QD�kAD{����	����ڐb�ǜF�&�L�A��\@d�r_���[�?���>(+�aG%�xSP���A	o�����ZX�I�7l�n�B�B����$����y�4�a`���o�y�[A|0�c5������dW��D�2Vi!0��c �R�
0p��Rɯ����|�3�un�CZ8�TDo0��@���y"���S���',�4���o���g`�����F'P�keq���t`�T�s�o*��sҸ��H8]����uy��v��=��� �$��duv��v2�v]������>7�f���W/w��N�8�%S����ډȻ$ʼ�i ������О4�]Sn#Ŀ�(S�' ��^ŝ��k�WS)2\�PE���/���Ae�#=� ^��;C��B�j��Q�)�z���/v �ܚ/�v��� �ѣ��]��W���Y��%s.�s����!������t�!g�Ĥ�>)$�f�z�T�p?\�H)��xQ��("�����	���5�ʀ���Jذ#�;ګ�`���&T!��������k3O�!���B!7ЂB5�!uzݢ��?`�_l�L����A�4D	��BW~A:�k��zz�>Fx����buz��$��P@?c/��H�eፄ۱� �6�g�Io���p����5��R$������C�&���E��F�JR���rC��b-%�����rN��T��E	�1�S!FCaǥj�x��*�Qp��%Ǚ���B��QթË��&e��d��cZrv�o�� �CK ��r�@}U����zv'vOMk��U��{��X���h���.��7��x�k��S��* ��@���Pgޙ:xWJU�6��-l����ˊ�����NR<�=�t�"1h�i�.�N8]�*n����+K5�D�J��]���#ͬl�-;L��ZE��`�J��M�O�s��nEV$����24�ѯ0^d�%PJ~�������!�$��%��"ɡ@�M:W��4�@;K��qp�x���c�Ǎ�$������I��a�� ���
&u+.#T�H��p��hd���2}��"us2�k�)�C��S�wW7# ;�=A��I��2��1�ԓ{�)ŷ�ظZ�f4�:�|����F`Ϻi�`e���<�i&�ʧ���I�+�p��M8!�0�M�� Λ�w�cR�٢x�q�Xy�g���d�m2���x��>���1�'ѷ��,'��siy����Ӹ�����5t�uB�����X����&c��{���h~6��T
$,�L#�RH8:�̤ɼ�A��#�CV:� ��^�
�j�Л���P��,�n�X�*Zy�0�\N����.%z��h�b?b��5���zǙD�dO�R�.��ԍ�#UDj/QHik�N�����7�T�,;����T���$l�az//����S�&��?�s���{P�*��aP>U�X�S�qh�찃s�£LR6ރ#inyP""��kJi磜��p�9�����v��$1����q��9��KN�8&�|�Q��-=��į49Q﷐p��T��#��td<=J�*�R%�ލ1�!I]�N�� ���ѧ8n����&D`��/E0��������;}�#�ץn,N1��;�@{�-����"DmJ1�r$O0��N}d&'�9�g��W���X�7XŶ�L���2�F!E��	:7Ά�Է�w�/S���ҟ`B��eL P������k�Ӳ��������TEL��žQ��;7����b���q�}ԅ��u_<�"�EW9��%�A���b$F��<�%�*���OLO/|�fxrjK��;�-�뎒.==2�W�� ���n4q�{�}�����
Z�ynV���о"�&ԥ�C�X$�SF,�N�mgյ�v��߱�b�X���&HS +��W����oǃ� ��U��Zg��V�j�������oK-�<����0V�r�[a\����`H�q�P�Y��)��Fک���K[�ƅ��p��J��ޠ��53�?J�i��MhP�����N9sS��q���-�r��(��ja��ץn��!�v���abw�{Ly���j떡(ԏ�k�7��'w�/��&�|g헴#�[������;�w�ɭ��x�����q�}�~f��Y[5E�N�I]��rhKE}M�z�_����+���0W�,�ǣ(w������wy�Z�Z�/u����Y�_�3����1s�"Ԙ��/�ՙs�I�:���^�o�>�=�o�W�7U��+!?�{�v{=MK�|���ѩ��䨹���C?��v|�)��P������}F��;��U��R��tf�s������e���\ ���i�|"�~P�V���}j�~V�WM�]~�����1C7����>��ަf?-�|�.�M�8ù��B��9��)���Q�>�A~Is�:���9�d����]�vQTV�z�\��5|<�� 0qw��~3:�$ɗU�e�;��u�>���7G����!.E��RRab�FL[pwW&nj�6�7��v��l�vq�T�KJ��;�����|�G�/�� �([6��h���I��mK1R�0N�W��x��u7�1 �}t�h"��[�8
@8�:̕�N��wd��i�����6_+q�������C�'<l0��!���$��q�0w�acRz*���0���n>zjY!_�)15ɟs㖔���$��pNwe*���L����vprl)�b�/�ۦ�7E`k������� �΂��DF��I2��K����k�%��|\��,�|�ilڹC�ə��� ��AIuw%E��������e7C���c�\!{ew�Z|2yӤPm�X�f:�~��љ�2���o�o�L˂��s�9���t#����Z�L�����L�\F���ڶ:�=S��'Yv�#���K�%r���S�� �M�E)2!46JLm���,`x�����1�����&��C�=Y��٤�[C�i{���C.G�X��N##�[���]�A�X���a�[_GoH뷹�����j(�C!�ȕ���Ɇ|W��z�{[�ɶ�H�M,� �O=̠��+���u1K�u�t��.��j�R�{;�)���md�	��n���(�l���j(�� ��E(�*ܵT�^�AB�;���=��|�N�$��__L��)N��>�1��[(�*z�d�	mmOsʹԗ�FX�@Z����bi��z�^!�����Ԃ��Pv�IuT)[����Z$w`������xlk�<��w�cZD
��WX�}�T͐ `c��!�����m v�uV�Dk��L灶գ͈�k�s�����P��:�	��Օz�����)�4qz���w˰�cEh�Z�ΌMvyuK`�
%��1�����IMn	TF!"`�SѝN�I�F�H��r_ͅ� !�H�Fná�˂#�a%�wl1pJHzY
f78Ó4XR���f#�(L�JuC!�;J�[u�JĺO�QN��Er7��s\��`D0�/l�AL�%A&�$��`�
�,gU��γ}+�v��fc�u2W�5�5�?� 1`i�^��yE�����(-He�j�s�ض�S��pX��k�W]M�
�eV���:
	.fhJV2hwq��B\���N}r�&N*��B�RL��fdp�]x7���&��n'�`��z�����$��QWU�s�����Y�P]�
i�z'���/\:�۩_�l��>~)�f,(�O�UcN�����8�$h6&�]3"�Lu*ºD~nh���uؼ��������Se�l��3�`F�F�blЉ����T�{#��w6
cf^O�A'��q ��ݍ�(�T��W�E���o�/7����E��ˣ�5ʚ#�8�<��I��ws��C�(_Y�gp�oͪ�WwoP3Uʴ��L��j��6�����:!����k93j��l�rCh��4+9 ����v]V0�{-I�<�r�t���ai![�<�?`�k`�.�#d�v�#��\�O��<
b����/��GX7�ˡU<l`	/���:%���X�0fG�t8hF�8�n�:z'�������>lȴ�C]#�嶴��`[&��TA��)	a�3뭲��\{c7A�2�퓕�� �܉�zSas��8T1&��Ц�;9���n�s��撹��T�fE�A�\J����쑻�̨����XڎC���꨽���=�F.B�]�v:�dϣ�Y}���p�*]�۪���v[���/�����m@N�����M�]�k1����9��1m�jFZM!�������-j�=V=��*w�ed֩�쵩���ؖ����6���x�Pdvk��(�nv���M��E
	6��q�2��@s�ho�3�He�R�� 6EvFJl����{�Q���ڡ��kL���_���m�9n�=�{@糐�{'-	�ƶ�0[3����D�ԭ���f������T[��d�N��n�M���쮻��A�J�Ӆ�o"����x;��nW�$.��Y�o��,��J	j׷5�7�ZX{�%�Njn���{^���.�؛Х�K�6�i:^�I���6Ig�Úu���J�׎�8 ��Դ������e8�f������f���?�,hvF��UMlm�r�Hz�]i�éR���8ٺ�.��q�@�&�8X�����~i�p�s�����x�zb�q��	k���=������3���l�.�wwQz%�{��Z���ܹ% IB�kr�	UW�O��2/����jA��%%���&F=\�2h�
W;��*��}BB�>2�j���q��p@� ���!��eH>�O��-v#�a��ڶ����.y[j�-	v����('��d�����$p��S\C��˛l��;A��ʽ�,A�r̄���Y�I�h�ҧ��J2��M��
���o��hO�#i�/$�Ӫ��;{������~Tq}�Zn'S ��Q��N��`�)�]��[�V|���䓶�l�<��Ħ��'��2m�e!�v��KM	}�"$��m\�s��Am�ձ���˾��v�H3�i��òk/��R� �	ĵ�C\�6�o�T%l�^t!�E�
����B����F���[6��=�C���I��W�I�����g�{o.�Z�`%��&��a��c����^_�H������5 {b`�F�0)��Hc^�uO���@�Ík���2o�mv9�%��h�J',��T�34)���f�M����۬��8z��&'��p����=��wA(ǯ1\6;�zXH�eieD��d�D��f��6�T��q5�MSТ7�x�F�D��O/���'QH�P2�I�{Y�2	�r{�̜�7�ʛR�g��sckz'����l��H�tdi�я9��7��ޣ�qc[��v�2q����Z���29��D���8�J����).G�ۦR(�=���3N(6�r�4ZN
/*k�U�06E/~X|�g]LN�Cj�ĆB�"^�p/B�!CĨ��B�TWj�v`N�c�H�vJRJ
f���\M@�B�Ld��O��oe�KU�R�O,R�ʙ�P�RXiM[Ѳ��� ���$� �`܂� ;S{M&46��Pt�u>��px�! ��@u�J2Ա<ʁ�Q���^W0�_|p�N������R�7���y}�c�!"���6	}2@�1aY��CiyaX�R�Pk���<:^�� ����87�1,W"	�d(��,�#r��膶���y]�S!=�'�^��X�Ӹ�X�d �7��O潸�R:��_΂��Ь��j�2�l����N7�^��� ��㕼��K_T�1�������'B�et`�
���0�CF��<"Vbq�?�����X`��j�in���S'e��қ��Unq犫�)��G�ʎc%n���i�
��Ti��%_����w��g�	�Q��S�(g�}��L�y!����&����X>�C�}<:>�G��D�&�U�>&�y�o�:)։vZ�C��/�������͌���԰S4w���>5�W&�@F�qz��}y�>�xa>��|P m(��K�c�P�EP>�<V�̓ʣ�p�}��D��K1���:����|�N��,��vF`����SN��V�PQ�-�PM/qս�O��׉S-mQ^�����0B��������H(�*�6sE��qm��L4Fg��_����N� ���M0]Q*�!��:O�h�kCg�_*�����[D`�V��q���,�+_�&:i,�\��%j����*t�YZ�-��FyB��i�G�)vN��UڦVVE���q	}�,����/�Q����%x������7���d�ηV�+����]n��(� آŋr��-���\�F���.���X[�np)V��i"v��K�����.�-͂����O���E� /l�  �
��d���r���pV�$������暊=�� ��N^ Do���*x����?����!	$��+5�r�������e�\�Mk��!V�����q�Fw��z1	$2� я8d��*
Q�`�U�W��ݜ��q?KI��((NQ�)4Yg�P.�Ef�k7�Hs��Ҵ7�2ew������W�����f�]V*�QE�"�(��:8�$&�dg	��'�檺:��_xz6靈?��b�7W�Ʈʷ;mk�-[	Bx�����ȶr���;��ӆs	x�[���FsKw�^����o�w1E�
��i����e���������I���|=!n��Є�4����^M�yӥ���mG����%z�W;6�\�j�
I���<��43I�'W
�Ӽ��:��!v��K���w��l���1�O:��*o�=�ʍ��Olr}��j�8}���<0n������7芭�R8��6��'?���u��1�T\x��ZKɸd��ϔJ�������<O�kgX�n�U�R�EG���ҟ6��ST��>��gQ���g	����C��+(��S�u��� 9-��5��vƪAW�σ����6��<U/�ԇ�6��[���<}��4�l�ۗy�i.�O��v[q|���5@W=��"H�ȴŕpy����=�|�J�)��,�*"��rsmݔ%�ٺ*|f==}�Cc��ݛ|rm���i��]\�k��BҤ��	r!h"�@��������f��r��٠\.�7ä�o,X���v:xQu!��|�<}m�8�ƨ��˕����6�v�f�Ŋ�k|�5��oɠ�Ѕzí��$��A0H��{Ao�h���%���>:&":���KW�@¯�l�{r0�����~��Uwh'A
IDX=6;4�O#*�|�z�q���i�.%�PO7���H�$?�6�,:M*-����Q� �M�_|�^:>KK��b�$�CwL�g\�޺�]q��E��ұ_j��Å��\j�(Ji�YT,A?��6Y �G�Ʃ�����g�勇��m�D9R	H1��Ԝ�t��j�u��χ9�Nrɡ�/K���Cd��tЁ�N��|���=�2�5&2���]�jfS�&P��\�D:��t����x�V����ޏ&7ְV@��Hx� �P;�ů�g�&�����8��B���^+f��8G�3�\[OD���wK8NW�ҾG�cf���{��g�b��F�Ӗn�*�7\O�&_�#�M�b�Wt���j��-��d�����a`�Y"�K�P�̾R���Ā���U������ឳ�91+�HD�)�̑)����qL_8��*�02���屶|4��
<ddB?$���\Dw;�]Td�-�I7�dR�[��u��)gF��@A!34���;O�}��S$�g���;���R!Jj�.c.Ro��$S4��C#F�J��N#X��)��z3P�(�]$+=����kl�d��.!\��3�D�K�|����$�-*��)�o�9�ƚn�*�Te��PZ�s��pn�/W1��!�"�[v�%O�X�Q!���dŷ'.��O_�@��ɞ4���S�m
�Iᗖ_�+�� ����{�O�fJĞ�� (�^��鱬�</��Xdz|L����|c�a"ߺ#�����<aN�yZ��V��p�P��'��s�a�BL,��d �GR6����ԥC��'�h�ľ҈��TㇶN�3Z����D��cӑ��zu���杧�S���rҪ�\��3u�u�8Mn".Qt<χ���>��C�[!t���*�[}�gr��F�`�k(��A��W���ԃ�pb��g����%�kr�4Kb����s�3����K�֭vI����1Ӻ��F1/ā�{z"���\�����E@��ƭ���QE��x�O�IOx�Iz��R������%4���)����K���o}=Nߨp�r�,�%%}%��,B�����u��}}e�g�[uu�P���.)���<˯��tM17�v��׮�]#$��8D$�i��ڢ�~���`��î��=���m����Yj��|Ҕ���a��Z�X����χ�'	^�M�}�ˡ�����D���c�5���#�>�0�u�-˜��t*���9h�U��h�'L���@�*0V�-VZ3o��)��\��a"U�8��A�.�3�YD�\w4Z�=	AT��b�����-�N|P*����oTl�i6/�X�xD�"ȋ�8�u���yY�⢼�)4��#�C�5��
EF&����*xr�����-ϸ��3W@����#V��qJ�#3u?dir^E�]��P��x�t]Z��n(��N�1�h�՘K�@�(ϓgx-��
bJ��G���)�!�U�%z�+f졁n[����{Q��mەr�%,�lتUش+';FA�7��۰LFT._,;�-�Wg�pGի���`��ƻ��]�M���L����vҚ�������-������ӥߡ�´��*+B.�vfߢ�`�2�lGy�VR����R{2Q�f�e٫d?VdU���&��s����oo���ո�ZM(4f�9�$kW(�N����P?t��s���e��za����ihK�'�fP��K�Л�kJslMљ�1=���2��d�����K�/��*��(�P��aU��,3Ś#���{E
�
ds����kV��$�\�1�BW�2����[x�@����vf��7��Y�p�����^��Q�<U6���� G��C�z��J&3�.�ݗ��
�f�bC�� n��^�$�*�-U��zx*����x]��Z�M�����juw�<n�MG�0�� �}���j�X=�d�qA�"��	Qb�d;��^Mn� H��6�B1�x̢� ���I�26�+����X�E�K��|Q��3E	�D&��L���r�2�UU�M��ʩ���}\�V�V�, ��R7eF77K��D�U7;�Ң���@^z:S��y�R�"���6� JMG�+a�N�Ұ[V5�x�f7L�z��V�_���P�W������g�������E���9z*�2O^Š���p�H��L�$͛��c�C������q�EA�yI�/=Y��(1�'��ov���O"w���eֵt��i���
������	�A1�� W�^��8��Yxa�}��|>@���w�)^!S�5v3��tZ��om�7˯��e���/x�g-��A|�,)t��@.��r�ձ�A
#�L��b�[���~���ji���RQ=�v*�X�����%�F�Z�m��W/�/|T�-	���Ŭ��>����E_�q!�jݱ/�ۇ��JR�z&lu���YB��k�2z��ߌBOi�q����0�/.��V�Q2�e�|TJ~�9� |����"]�L0g)��LC�龐��2�G�0�b_l��_E!`ޯp}w�j���9��cP��Wo���QH���:���ŉ��Y�o�˸6��G:hn��BG0R��xW,�H��y�@=�c|�.ڟ��>hc�Pbt��WYI`�qHpI�➇;�&�x����c���ړ�d��v��K��eH�(B�=6clDYB`��(?c!h�ߝ�C�=�
�nv�����.]����u��$����*���̋[�#y���KF�
	d����� C��� a����}���wlz�p���~7�8��f�X��*�oH���"AG��E���Di��s6���a38ۻ4�G��	��ɥ��9]=����j�z746���;>N$�y8����[�	/�^��O�5x���$x[�=��o���õ��֥�`��_̹�V�s�!�nH=��=1�`�Pe�=b��&BZ��*�8G+Z��� ���8��r���:����{����@:M���>E�o��S��0�7�����;.�H{rp�ɾ�2��Q�5n��^��fz$74�2�<\�