U�Q�e�E�M���  ���E�E��]���������������U����E�E��M�Q�UR�EPQ�e�M�U�Q�e�E�M��  ���E�E��]���������������U��j�h'^' d�    Pd�%    Q�E�    �EP�MQ�UR�	  ���E����E��E�M�d�    ��]���U��j�h�]' d�    Pd�%    Q�E�    �EP�MQ�UR�/	  ���E����E��E�M�d�    ��]���U��j�h�]' d�    Pd�%    Q�E�    �EP�MQ�UR�O	  ���E����E��E�M�d�    ��]���U��j�h�k' d�    Pd�%    ��h�M��E�� �3( �E�    �M���3( �E�   �U��|�+ �E����EȋM��@   j@�� ���E̋UȋẺB�E��M����M��U��@   j@�� ���EċE��MĉH�E��U����U�jj@�M���� �E��E�� \8( �E��M��d9( �M��Z�
 �E��}@w�U��B�E��MQ�UR�E�P趥 ���yjj@�M��� �E��E�\8( �E��E�d9( �M���
 �E��MЉM��E�	�U��U��E��H�M��UR�EP�M�Q�U���M��P�E�
�E��E��M��O/���E   �M��Q�U��@   +EPj �M�MQ�� ���E�    �	�U����U��}�@sH�E��H�M��U��B�E��M�M����\�E�E���M��Q�U��E�E��E��M����6�E��멋M���  �E������E��M�d�    ��]� ���U��Q�M��EP�MQ�M����U��B�P��]� ������������U��j�h�7' d�    Pd�%    �� �M��E�   j��� ���E�E�E��E�    �M��M�U�R�Mԃ��EԋP�R�EԋH�M�j@�U�R�Mԃ��EԋP�R�E��E�j�M�Q�Mԃ��UԋB�P�MQ�UR�Mԃ��EԋP�R�M���  �E������E�Pj �M�Q�j� ���U��U؋E�P蛷 ���M�d�    ��]� �����U����E�����E��E�    �	�M����M��U�;U�s�E��M��R�U(�����M��U���ҋ�]����U���0�MԋE�P�MQQ�e�U�E�Q�e��M��U��b  ���EЋEЋ�]� ���U���0�MԋE�P�MQQ�e�U�E�Q�e��M��U��b  ���EЋEЋ�]� ���U���T�E�E��M��M�U�E��M��M�U�E��M��M��U��E��M�+M����A�����B��t5�M����M��U����U��E��E��M��M��, Rj �E�P�M��ͷ��뱋M�U���E��]�������������U���T�E�E��M��M�U�E��M��M�U�E��M��M��U��E��M�+M����A�����B��t �M���H�M��U���H�U��E�P�M��"  �ƋM�U���E��]��U���4�E�E��M̉M�U�E��MЉM�U�E��MԉM��U��E��M�+M����A�����B��t8�MЃ��MЋŨ��ŰEЉE܋M̉M؋U؋E܋�
�U؋E�f�Hf�J뮋U�Ẻ�E��]����������U���0�MԋE�P�MQQ�e�U�E�Q�e��M��U��	  ���EЋEЋ�]� ���U���	�E���E�M+M���A�����B��t�MQ�M�\  ��]���������U���,�E�E��MԉM�U�E��M؉M�U�E��M܉M��U��E��M�+M����A�����B��t �M؃��M؋Uԃ��UԋE�P�M���  �ƋM�Uԉ�E��]��U���0�MԋE�P�MQQ�e�U�E�Q�e��M��U���v ���EЋEЋ�]� ���U��Q�M��M���k���E����t�M�Q�j� ���E���]� ��U���`�M��, Pj �MQ�M������U��Ef�Hf�J�U��E�H �J �, Rj �E��$P�M���$�δ���M��U�B@�A@�M��U�BD�AD�E���]� �������������U��Q�M��M���)���E����t�M�Q躞 ���E���]� ��U��j�hk' d�    Pd�%    ��(�M��E�    �E������Ẽ��E��E�   �E������MЃ����  �M�d�    ��]�����U��j�h�]' d�    Pd�%    Q�E�    �E� 4, �M�A �E�   �U���+ �E�M�H�U�E�B�E� �M����M��E�M�d�    ��]�U��j�ho]' d�    Pd�%    Q�E�    �E� 4, �M�A �E�   �U�p�+ �E�M�H�U�E�B�E� �M����M��E�M�d�    ��]�U��j�h?]' d�    Pd�%    Q�E�    �E� 4, �M�A �E�   �U���+ �E�M�H�U�E�B�E� �M����M��E�M�d�    ��]�U��j�h��' d�    Pd�%    �� �MԋEP�M�薒 �E�    �M�Q�M���v �UԉU��E������M��� �E�M�d�    ��]� �����������U��j�h ]' d�    Pd�%    Q��SVW�e��E�E��E�    ��M���M�U���U�E+E���@�����A�х�t?�E�E�M�M�}� t$�U�E�
��J�H�J�H�R�P�E�E���E�    ���	�M���M�U�;Ut��j j ��� �E������E�M�d�    _^[��]����������U����M��E��H�M�j@�U�R�M����E��P�R��]������U����E�E��M�Q�UR�EPQ�e�M�U�Q�e�E�M��;  ���E�E��]���������������U��Q��E���E�M���M�U+U���B�����@�ȅ�t �U�U��E�M����E�M�f�Qf�P봋E��]��������U��j�hQ~' d�    Pd�%    Q��LSVW�e��E�E��E�    ��M���M�U���U�} vJ�E�E��E��}� t'j �M����	 �, Qj �UR�M������E�E���E�    �M��M��E� ��=�	�U���U�E�;Et!j�M���	 3Ƀ���t�U�R�� ����j j �� �E������M�d�    _^[��]�������U��j�h�' d�    Pd�%    Q��TSVW�e��E�E��E�    ��M���M�U��H�U�} v4�E�E��E��}� t�MQ�M�������E���E�    �U��U��E� ��*�	�E��H�E�M�;Mt�U�R��  ����j j �?� �E������M�d�    _^[��]����������������U��j�h�V' d�    Pd�%    Q��SVW�e��E�E��E�    ��M���M�U���U�} v-�E�E�}� t�M��A�M��A�U�U���E�    ���	�E���E�M�;Mt��j j �� �E������M�d�    _^[��]���U��j�h!�' d�    Pd�%    Q��SVW�e��E�E��E�    ��M���M�U���U�} v4�E�E��E��}� t�MQ�M�軍 �E���E�    �U��U��E� ��;�	�E���E�M�;Mt�M��� 3҃���t�E�P谗 ����j j �� �E������M�d�    _^[��]���������������U����	�E���E�M;Mt!j�M���	 3҃���t�EP�G� ���΋�]���U����E�E��M�Q�UR�EPQ�e�M�U�Q�e�E�M��  ���E�E��]���������������U����E�E��M�Q�UR�EPQ�e�M�U�Q�e�E�M��Ks ���E�E��]���������������U��j�h��' d�    Pd�%    Q��xSVW�e���x����E�E��E�    ��M��U�E+E���@�����A�х�t�E��P�MQ��x�����������Q��U��E�M�+M���A�����B��t$�M�M�U�B�E�M�Q�U�R��x����ק �j j ��� �E������M�d�    _^[��]� ��U��j�h�7' d�    Pd�%    Q��SVW�e��E�E��E�    ��M���M�U���U�} v'�E�E�}� t�M��E��M�M���E�    ����	�U���U�E�;Et��j j �8� �E������M�d�    _^[��]���������U��j�hq�' d�    Pd�%    Q��XSVW�e��E�E��E�    ��M��H�M�U��H�U�E+E���@�����A�х�t:�E�E��M�M��E��}� t�U�R�M�������E���E�    �E��E��E� ��*�	�M��H�M�U�;Ut�E�P��  ����j j �U� �E������E�M�d�    _^[��]���U��j�h]' d�    Pd�%    Q��SVW�e��E�E��E�    ��M���M�U���U�E+E���@�����A�х�t3�E�E�M�M�}� t�U��J�U��J�E�E���E�    ���	�M���M�U�;Ut��j j �� �E������E�M�d�    _^[��]������U��j�hQ�' d�    Pd�%    Q��PSVW�e��E�E��E�    ��M���M�U���U�E+E���@�����A�х�tP�E�E��M�M��E��}� t'j �M��c�	 �, Rj �E�P�M�莨���M�M���E�    �U��U��E� ��=�	�E���E�M�;Mt!j�M���	 3҃���t�E�P�~� ����j j �|� �E������E�M�d�    _^[��]����������U��j�h�\' d�    Pd�%    Q��SVW�e��E�E��E�    ��M���M�U���U�E+E���@�����A�х�t-�E�E�M�M�}� t�U��M��U�U���E�    ���	�E���E�M�;Mt��j j �� �E������E�M�d�    _^[��]������������U��M�]��3�����t�MQ�_� ��]��������������̃��X� �������̃��x� ��������+I��� ��������+I����� �����+I����z�������+I����u{������̃���� �������̃��� �������̃���� �������̃���� ��������+I��H� ��������+I��8z����������+I��{����������+I��(����������+I��� ��������+I������������U���$�M܋M���   �E܃8 u� h�  hL�+ h�+ h��+ �Þ ���6� �M܃y( u�U܃z$ u� h�  hL�+ h��+ h��+ 菞 ���� �E܋H$�M��U܋B�E�M�M�U����E�E�M�M��U��z t�E��8 v�M��y u�U��z u� h�  hL�+ h��+ h��+ �� ��葥 �E�� ��]��������U����M��E����E��M��y u	�E�    ��U��E��J+H���M�U����U��E��x u	�E�    ��M��U��A+B���E�M�;M�u� h�  hL�+ h4�+ h�+ 聝 ���� �U����U�E�x u	�E�    ��M�U�A+B���E�M��Q$;U�s� h�  hL�+ h��+ h��+ �'� ��蒡 �E��H$���U�9J(w� h�  hL�+ hH�+ h�+ ��� ���_� ��]���U��Qf�E� f�E�  j�E�Ph�   h��  �MQ�`( ��]���U���0�} t�E�8 t�} t�M�;Uw� h�  hT�+ h�+ h��+ �x� ���� �E�M;Mvjh��+ �M�����hԠ- �U�R�� �E��M��U�E�M��E���]�����U���,�} t�E�8 t�} t�M�;Uw� h%  hT�+ h�+ h��+ �� ���[� �E���;Mvjh��+ �M��^���hԠ- �U�R�� f�EP�d( �������   �U���   ;�u'f�EP�d( �ȁ��   �U�����   ;�u�h2  hT�+ h(�+ �W� ���� �E��%�   �M���E����U�
�E%�   �M���E����U�
��]���������U���D�M��M�������E��8u� h7  hL�+ h�+ h��+ �Ӛ ���F� �M��Q$�U��E��H�M�U�U�E��M���U�E�x u.�M��Q$�UЋE��H�MԋUԉU܋EЋM܍��U؋E؃8 u� h=  hL�+ hp�+ hD�+ �X� ���ˡ �M��Q$�U��E��H�MċUĉŰE����M�ȉMȋUȉU��E��M��P;Qu&�E��HM�U�;Js�E��H�U�
�E�9Hw� hC  hL�+ h`�+ hH�+ �ؙ ���K� �M��AE��]� �����������U���D�M��M������E��8 t(�M��9t h  hL�+ h�+ h��+ �}� ���� �U��B$�E��M��Q�U�E�E�M��U�ʉE�M�y u.�U��B$�EЋM��Q�UԋEԉE܋MЋU܍ʉE؋M؃9 u� h$  hL�+ hp�+ hD�+ �� ���u� �U��   j�M���- �E��H$�M��U��B�EċMĉM̋U����E�EȋMȉM��U��E��J+H����]����U���,�} t�} t
�E;Ew� hD  hT�+ h��+ h��+ �r� ���� �M;Mtjht�+ �M�����hԠ- �U�R�� ��]������������U���,�} t�E�8 t�} t�M�;Uw� h  hT�+ h0�+ h�+ ��� ���k� �} t� h  hT�+ h �+ h��+ �З ���C� �E�M;Mvjh��+ �M��F���hԠ- �U�R� � �EP�M�R�EP��� ���M�U�E���]��U���0�} t�E�8 t�} t�M�;Uw� h2  hT�+ h0�+ h�+ �8� ��諞 �E�M;Mvjh��+ �M�讷��hԠ- �U�R�h� �E��M��U�E�M��E���]�����U���t�M��M�������E��8t8�M��9t0�U��:	t(�E��8
t h|  hL�+ h��+ h��+ 蝖 ���� �M��Q(�U��E��H�M��U��U��E����M�ȉM��U��U��E��x ��   �M��y ��   �U��E��J;H��   �U��z0 u2�E��H(�M��U��B�E��M��M��U��E��ЉM��U��E��J;HuT�U��z0 tI�E��x4 tB�M��U��A;B4w4�M��Q(�U��E��H�M��U��U��E��M����U��E��M��P;Q4u� h�  hL�+ h��+ h��+ 薕 ���	� �E��HM�U�;Jvjh��+ �M�����hԠ- �E�P��� �M��
   �U��B�E��M��QU�E��P�E���]� U���t�M��M������E��8t8�M��9t0�U��:	t(�E��8
t h�  hL�+ h��+ h��+ �� ���`� �} t� h�  hL�+ h �+ h��+ �Ŕ ���8� �M��Q(�U��E��H�M��U��U��E����M�ȉM��U��U��E��x ��   �M��y ��   �U��E��J;H��   �U��z0 u2�E��H(�M��U��B�E��M��M��U��E��ЉM��U��E��J;HuT�U��z0 tI�E��x4 tB�M��U��A;B4w4�M��Q(�U��E��H�M��U��U��E��M����U��E��M��P;Q4u� h�  hL�+ h��+ h��+ 输 ���1� �E�� 
   �M��Q���E�;Pvjhx�+ �M��'���hԠ- �M�Q��� �U���U��E����E��M��Q�E��
��U��B���M��A�U����U��E��H�U����M��Q���E��P�Mf�R�d( ����%�   �M����   ;�u+�Ef�Q�d( �Ё��   �E������   ;�u�h�  hL�+ h��+ �ƒ ���z� ��]� ��U���D�M��M������E��8t8�M��9t0�U��:	t(�E��8
t hD  hL�+ h��+ h��+ �m� ����� �M��Q(�U��E��H�M�U�U�E����M�ȉM�U�U��E��x ��   �M��y ��   �U��E��J;H��   �U��z0 u2�E��H(�MЋU��B�EԋMԉM܋UЋE܍ЉM؋U��E؋J;HuT�U��z0 tI�E��x4 tB�M��U��A;B4w4�M��Q(�U��E��H�MċUĉŰE��M̍��UȋEȋM��P;Q4u� hW  hL�+ h��+ h��+ �f� ���٘ �E�� 
   �M��A��]������U���H�M��M��/����E��8 t(�M��9t h�  hL�+ h�+ h��+ �� ��耘 �U��B$�E܋M��Q�U��E��E�M܋U�ʉE�M�y u.�U��B$�E̋M��Q�UЋEЉE؋M̋U؍ʉEԋMԃ9 u� h  hL�+ hp�+ hD�+ 蒐 ���� �U��   �EP�M��b% �M��Q$�U��E��H�M��U��UȋE����M�ȉMċUĉU��E��H�M��U��BE�M��A�E���]� ��U���D�M��M������E��8 t(�M��9t h>  hL�+ h�+ h��+ �� ���`� �U��B$�E��M��Q�U�E�E�M��U�ʉE�M�y u.�U��B$�EЋM��Q�UԋEԉE܋MЋU܍ʉE؋M؃9 u� hD  hL�+ hp�+ hD�+ �r� ���� �U��   j�M��D$ f�EP�d( �������   �U���   ;�u'f�EP�d( �ȁ��   �U�����   ;�u�hR  hL�+ h(�+ ��� ��謓 �E��H$�M��U��B�EċMĉM̋U����E�EȋMȉM��U�����   �E��H��U��B���M��A�U���   �E��H��U��B���M��A��]� ���U���D�M��M��_����E��8 t(�M��9t h�  hL�+ h�+ h��+ �=� ��谕 �} t� h�  hL�+ h��+ h��+ �� ��舕 �U��B$�E��M��Q�U�E�E�M��U�ʉE�M�y u.�U��B$�EЋM��Q�UԋEԉE܋MЋU܍ʉE؋M؃9 u� h�  hL�+ hp�+ hD�+ 蚍 ���� �U��   �EP�M��j" �M��Q$�U��E��H�MċUĉŰE����M�ȉMȋUȉU��EP�MQ�U��BP�~ ���M��QU�E��P��]� ���������������U���p�M��M�������E��8t8�M��9t0�U��:	t(�E��8
t hA  hL�+ h��+ h��+ �͌ ���@� �} t� hB  hL�+ h �+ h��+ 襌 ���� �M��Q(�U��E��H�M��U��U��E����M�ȉM��U��U��E��x ��   �M��y ��   �U��E��J;H��   �U��z0 u2�E��H(�M��U��B�E��M��M��U��E��ЉM��U��E��J;HuT�U��z0 tI�E��x4 tB�M��U��A;B4w4�M��Q(�U��E��H�M��U��U��E��M����U��E��M��P;Q4u� hU  hL�+ h��+ h��+ 螋 ���� �E��HM�U�;Jvjh��+ �M�����hԠ- �E�P��� �M��
   �UR�E��HQ�UR�| ���E��HM�U��J��]� �������������U���P�M��M������E��8 t(�M��9t h�  hL�+ h�+ h��+ �� ���`� �U�B�E�}���  w� h�  hL�+ h|�+ hh�+ 蹊 ���,� �M��Q$�U؋E��H�M܋U܉U�E؋M���U��E��x u.�M��Q$�UȋE��H�M̋ỦUԋEȋMԍ��UЋEЃ8 u� h�  hL�+ hp�+ hD�+ �>� ��豑 �M��   �U�B�E�f�M�f�M��U���R�M��� f�E�P�d( �������   �U����   ;�u'f�E�P�d( �ȁ��   �U������   ;�u�h�  hL�+ h��+ 證 ���a� �E��H$�M��U��B�E��M��M��U����E�E��M��M��   ��t�h�  hL�+ h��+ �[� ���� �E���%�   �M��Q��E��H���U��J�E�%�   �M��Q��E��H���U��Jj �E�P�M��QR�M��,  �E��M�A�U��B��]� ��������������U���t�M��M������E��8t8�M��9t0�U��:	t(�E��8
t h�  hL�+ h��+ h��+ 荈 ��� � �} t� h�  hL�+ h �+ h��+ �e� ���؏ �M��Q(�U��E��H�M��U��U��E����M�ȉM��U��U��E��x ��   �M��y ��   �U��E��J;H��   �U��z0 u2�E��H(�M��U��B�E��M��M��U��E��ЉM��U��E��J;HuT�U��z0 tI�E��x4 tB�M��U��A;B4w4�M��Q(�U��E��H�M��U��U��E��M����U��E��M��P;Q4u� h�  hL�+ h��+ h��+ �^� ���ю �E�� 
   �M��Q���E�;Pvjhh�+ �M��ǧ��hԠ- �M�Q�� �U���U��E����E��M��Q�E��
��U��B���M��A�U����U��E��H�U����M��Q���E��P�M����M��U��B�M����E��H���U��J�E����E��M��Q�E��
��U��B���M��A�U�P�h( ��%�   �M����   ;�uq�E�Q�h( ��%�   �U�
�����   ;�uK�U�P�h( ��%�   �M������   ;�u%�E�Q�h( %�   �U�
�����   ;�u�h�  hL�+ h@�+ �ۅ ��菊 ��]� �������U����   ��<�����<���������<����8
u� h�  hL�+ h$�+ h�+ 臅 ����� ��<����Q(�U���<����H�M��U��U��E����M�ȉM��U��U��E��x ��   �M��y ��   �U��E��J;H��   ��<����z0 u8��<����H(�M���<����B�E��M��M��U��E��ЉM��U��E��J;Huf��<����z0 tX��<����x4 tN�M���<����A;B4w=��<����Q(�U���<����H�M��U��U��E��M����U��E���<����P;Q4u� h�  hL�+ h��+ h��+ �_� ���ҋ �E��M��P;Qtjh��+ �M��Ԥ��hԠ- �E�P�� ��<����y0 uF��<�����<����J(;H$u� h�  hL�+ h��+ h��+ �� ���e� ��<�����   �   ��<����z( u��<����x$ u� h�  hL�+ h��+ h\�+ 訃 ���� ��<����y4 t)�U���<����J;H4w�U��B�M���<���9B4w� h�  hL�+ h��+ h��+ �S� ���Ɗ �E���<����P;Q4u��<����)   ���<����    ��<���������]�������������U���\�M��M�������E��     �M��A$    �U��B(    �E��@,    �M��Q$�U�E��H�M�U�U��E����M�ȉM�U��B    �E��H$�MԋU��B�E؋M؉M��U����E�E܋M��A    �U��B$�EċM��Q�UȋEȉEЋMċUЍʉE̋M��A    �U��B$�E��M��Q�U��E��E��M��U��ʉE��M��    �U��B0    �E��@4    �M��������]��������������U���p�M��M�������E��8t8�M��9t0�U��:	t(�E��8
t hi  hL�+ h��+ h��+ 蝁 ���� �} t� hj  hL�+ h �+ h��+ �u� ���� �M��Q(�U��E��H�M��U��U��E����M�ȉM��U��U��E��x ��   �M��y ��   �U��E��J;H��   �U��z0 u2�E��H(�M��U��B�E��M��M��U��E��ЉM��U��E��J;HuT�U��z0 tI�E��x4 tB�M��U��A;B4w4�M��Q(�U��E��H�M��U��U��E��M����U��E��M��P;Q4u� h}  hL�+ h��+ h��+ �n� ���� �E�� 
   �M��Q���E�;Pvjht�+ �M��נ��hԠ- �M�Q�� �U��B�M���E��H���U��J��]� �������U���D�M��M�������E��H$�MЋU��B�EԋMԉM܋U����E�E؋M؉M��U��B$�E��M��Q�UċEĉE̋M��U̍ʉEȋMȉM��U��:�!  �E��x0 t� h  hL�+ hT�+ hT�+ �p ���� �M��y t4�U��: v,�E��x4 t#�M��U��A;B4w�M��Q�E��M�9Q4w� h  hL�+ hX�+ h,�+ � ��膆 �U��z t=�E��8 v5�M��y t,�U��E��J;Hu�U��E��J;Hw�U��E��J;H4w� h$  hL�+ h �+ h��+ �~ ��� � �U��E��J4+H�M�U+U�U��}� ��   �E��H�U�
�E�+H4�M�M�;M�r%�U��E��H4�J�U��B0    �E��@4    �   �M�Q�U��BP�M��QR�� ���E��M��Q�P�E��HM�U��J�E��@0    �M��A4    �U��B    �E��     �M�Q�M��� �U��E��H�J�U��E��H�J�U��E���M��   ���   �U��E��H�J�U��E��M��A0    �U��B4    �E��    2��   �M��9 t(�U��:t hv  hL�+ h��+ ht�+ �J} ��轄 �E��x u�M��9 u�U��z u�E��x u� h|  hL�+ h�+ h��+ �} ���x� �MQ�M��� �U��E��H�J�U��E��M��   ���]� ������U���D�M��M������E��8 t(�M��9t ha  hL�+ h�+ h��+ �| ��� � �U��B$�E��M��Q�U�E�E�M��U�ʉE�M�y u.�U��B$�EЋM��Q�UԋEԉE܋MЋU܍ʉE؋M؃9 u� hg  hL�+ hp�+ hD�+ �| ��腃 �U��   j�M��� �EP�h( ��%�   �M���   ;�ue�UR�h( ��%�   �M�����   ;�uC�UR�h( ��%�   �M�����   ;�u!�UR�h( %�   �M�����   ;�u�ht  hL�+ h�+ �`{ ���� �U��B$�E��M��Q�UċEĉE̋M����U�щUȋEȉE��M�����   �U��B��M��Q���E��P�M�����   �U��B��M��Q���E��P�M�����   �U��B��M��Q���E��P�M���   �U��B��M��Q���E��P��]� �������U���D�M��M������E��8 t(�M��9t h%  hL�+ h�+ h��+ �]z ���Ё �U��B$�E��M��Q�U�E�E�M��U�ʉE�M�y u.�U��B$�EЋM��Q�UԋEԉE܋MЋU܍ʉE؋M؃9 u� h+  hL�+ hp�+ hD�+ ��y ���U� �U��   j�M�� �E��H$�M��U��B�EċMĉM̋U����E�EȋMȉM��U��B�M��U��B���M��A��]� �����U��j�hF�' d�    Pd�%    Q��`SVW�e��M��E�   �E��M��8����E��H�M؋U؉U�E��H�MԋUԉU��	�E���E�M�+M����A�����B��t�M�QR�n ���E��@    ����ދ ��E�   �E� �M����L   �E������M����z�  �M�d�    _^[��]����������U���$�M܋M��   ��]������������U���$�M܋E܃x tf�M܋Q�U�E܋H�M�U�U�E�E��M��M��U��U��	�E����E��M�;M�t��U܋E܋J+H���M�U܋B�E��M�Q�Wi ���U��B    �E��@    �M��A    ��]�������U��j�h�' d�    Pd�%    ���   �����������     ��������M�j �M��j� �E�    ��������U�j �M��< �E�������@$    ������A(    ������B,    ������@0    ������A4    �} v� h�  hL�+ h��+ h��+ �w ���~ �E�    �E�    �E�    �E�    ���ԋE���M��J�E��B�M��J�UR��������  �E�P�M�Q�UR��������  ����������} �  ǅX���    ������H��\�����\�����d�����X�������d���ȉ�`�����`�����T����EP��n ����T����AǅD���    ������B��H�����H�����P�����D�������P����L�����L����y u,jh��+ �M��C����E��E��, �E�hԠ- �U�R�� ǅ$���    ������H��(�����(�����0�����$�������0���ȉ�,�����,����E�������d����E�����������M�d�    ��]� �������U��j�h��' d�    Pd�%    ��   ��`���j �M���	 h, �i ��Ph, �M�跔���E�    �E�P�M��p���E��E�X/( �E� hT�- �M�Q�/� �M�d�    ��]����������U���   ��p�����p����x uǅl���    ���p�����p����A+B����l�����l���;Msi��p����z uǅh���    ���p�����p����P+Q����h����EP�M+�h���QQ�e䋕p����B�E�M�U���p����   �   ��p����x uǅd���    ���p�����p����A+B����d����M;�d���sSQ�e܋�p����B�E��M܋U����p����H�M؋U؉U�Q�eЋE���M�ȉMԋUЋEԉ�M�Q��p����	  ��]� ���U��j�hP�' d�    Pd�%    Q��L  SVW�e��������E��M��P�U�H�M�P�U싅�����x uǅ����    ��������������A+B���������������M܃} u��  �E�����}� v�U��������
ǅ����   �������x uǅ����    ��������������A+B��������������+�����;Ms�������#����O  �������z uǅ����    ��������������P+Q��������������E9E���  ǅ8��������8��� v��8����������
ǅ����   �U��ꋅ����+�;E�sǅ����    ��M���U�щ������������E܋������y uǅ����    ��������������J+H��������������U9U�s?�������x uǅ����    �����