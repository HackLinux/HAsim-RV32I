T���<����{�%4 �CK�]{xU��W��$v�tx���a��7q� :۝t�;�(�eȪ0�aI$�AS{�#����U�����Qv��G��Jb�Ft��TO>]
��[U]Տ������[��{����W�kI�%צ�@��j�W��Y���OR���d��y��ѳ
:Ԋ�C�wk��[�[�RF�&��Ԅ�Ԅ���	���Za��T�J+��vƭp�[}#F�ǐ��"���B��U���
�JPz��7��G�APoG��9��Z��K���pƽ�.	�SpŹq��̛v2h:E�ÿ��z�J7z�,,���h��[lP\Z�G��#�bo'Ldp�l �):�_�$w�,c� {}؂p�^�G�H���� �'M"HA���Fj�ʅ�|��l��WN p�&Щ=(�t�i݉�Z��,�`����4_��GA�-dWT����bPM�=V��r~`������'xl*���������h3�<ƃ1���a)�E��+	b!���I�R8�}�p.[(ĖXyT���Y���*i��D�<�}.�V6������XG{I�Ƅ3�S��;�
�%d�^�#JyE��3�=X}��[&+���b�h�6g=��E[�_ҿ�����9�W;�7c�T~��e+�#�:b�-��)Z's�M*Fe~6D���!�~G:,��#�ZA*��Jfb�3�'z�A`e�t�C|���4m�{��a��+_����%>٫���E��	���r��R�~k�8�VJ�t�q��v���s�8(�w����+��Ȓ����p#.��=ĭ���g�oK��|ݰs���Ź�X�ؿC#��Ng�"9�A�x>�H��Ć=��Z��]O��s��,�=��&�k>ON�x���n½~�@Ѭ̝z4���#E���.n���X�Ű��q5�QP����%u�� �K�3	��EL*J?���;��};�3�O�s����Р����E��r���a�y���hЖ�JOP1��q�ё���*�2ૈ4��'� �u��~q����#��Ǯ�Z7���/S�lN�&bp_Z#�$�!#���V$U�Ir`gZ+z���U�;��ޭs�i L�u�����]J�S K������Bf�p�5�
Q��Ʒ���3�V�ض�y��R9�׷�ɤo5��D<+���}�j�}��t
��Ϭ٢ξ�m��?ճf�a�5%@�t�r()y,h$�nFjA�%�9��o�7�.�?�����UT?��,r��Hi5�gcY�ǅe���W� �0{|�I	ڷ�wf�t i�5��(9y�^��r��q����%�\"�* /��0��46�!�m|�!���Z<5�*l�e�G�p�1&%��6�E�LF�N�~�[�E&S�)�r>a���Tn��e��w,�������������?�_������;�彭�q�5��?CQ?�Dٰ�l���E2�F3��,$GH]��^�:L���j�o#�{�6]�2�>�t�2KQd����;�*��d���v�~{��҅����K��{n���g��@�/쪡w��+�1��qKc]8n��6?8O+�9)a�dXw����.2S��m��R~�~C7�����nO�[�� �Ȃ��L������@��>���������x�l'E_���_&j��M��:aհ�^֗L�r��Y����cx��36��1�,�<^�e���SŹzk�bߌ���i�ĳ��$�*I�=Ì���ޞ!�5��PEws��w�*��U5��7�W�&�ghr�����*N��Q
6T�{���OgS��C׫)���}k'�@�u�~1���� ���U9$�ژ�")ނ���[BF�_����a�,�t�V@����	W'W�F8�)��r�4�MLYK�>;����u�x�J�X#�Fv���0��K�b�t�YI���(&��	����Bh�޲��a���[�5O�l,lc:\3�����2j~؝�K;�!
d���П�͸��v])�:��S.M~��^��Z(�^ JƷ����s����fOC��o��w�����1\���O�$}Yg�V�/�2"�?�ũ??qe�ϭԟ��I�WN
e7Նw������J�ݡD�5�:�&������_����� F}�^UɃ�����Q���{F3���贰II���ڟ��_Pܣ]����B�"���3��gğ����3��)Woc������?����U�~�y*�'T��3�o�]��G e�X 0��!H�=�I59�o�~T��K�3���'m���1~Z�Pq�LYq?��-�ߩ��l`�U�ip����oP\c!,U�����\n>�^��+�o����G���T��dM���}��tЦ�Nij��F������k-����`y��vqm̂l�W��b��*���J��>�,���I�'>O��6͠(5��P�&�����2Y)m��� x�ޟk%�Gp.�����)��!v*��I=���+����%Pa�f�wZ�`o_iU�� �'��^�����S���|[d64�u��raq!��pD�b��|�.ŀj�AX+��jk���FB��F�	�ïp��M��AD�\�Vb�G�J?��:! �r�Z8{f�\��Ѭ�Hܭ{���}$������yG�z,PKƄ@ȇ�"�ɨւ�6�%=4K���@gi�zG��iJ�t(,�X��M����þ���W�͑iD��`���;lNU_���
��q1O}�Q��r���@��v�����/6�Y�����aJI�)��SF����Pv��Fxr�Iμ����I�'{3��� ۣ�P���z���8�۩��C�~��0RR��HO:xR�z|r��Or��Gp��l7�DF4��FZ��d��i��&ݸj��;hDs��PI�~�x�;#�N�G:U<�q}����\8v������k���r�W�w�7|K�i����Y��n���xĿ�?j�O���T_����%Q����94��]�ûyyo�D���
E4�Z3�0�s~J~V�/�vvp�l�����m������;��F����/�R����c}A��'Uo����y�e�Jfd��G��-���Z��$
�	ܟ�2����'~(��J����H���&\����L��Λ�H��$z{�������&�2�WmlO���h��2�֢k@�\?�۷���JL��*��X��/�Ӣ�%�>�imV�zR�,�h6c�|A-�'����/����ǋ7�5f�C.|(�u���)�~��>=��s�J�(�5��vq�E��@3ESlS�`쟛��b�����.��Z�6��TO������S�pQ<��d<�h[�2|P<��,��EOrT��h�m�����]��J�?�����K:�XN<��;�v�!�Xz��^i��e$�pZ��г"=!#��K�gCz��􎟿Dz���H��K����<�U��7|1��`T�c@��]L���8?��s`����bg�	����.�_7� V
C�z�*�bZ<Z'�6�,��+%(z>1���KI��|%u�wly��[J1ּ.�["z��^w���P8m�дn����o�"����C���*@S�gs��������:�g�� �0�Z�'GD�󢠼�*�<�Zz�c-�����ǳ��oVv$�]�=�W3���&zm�RAʫ��y��La����̮��o��R���`��:�3G���!��1���N7- up�Xnhy�ǆj"7E+�[}Q���ޞ�	ka�uχ��ZP���t�H�����8ܚ�]	y	xb���R>v+��a8b���J������0
��/W�}e;�-�f_Y��,��Tjs:!�ܕ�G���-��o��������"ScY���˚��(��X̀��57�ؾ%��?,l�}k�#z,���)��Sȁs�p��b���������D|�=�Cc��s�>x�Jz�l�������g�[O5۷�:��V�U��N�V9�lJ�J��v	Ѷo�=f�9�E:�Q��$�VO�)O�I~LߍGX,�i[吞�JkȽ�DC\������L��s�6���' }衧l_�1Kr3��-fK.6�Z`�`-E�!_� ��!7��1jh��6�j�g7���,�7�j'�c��Q�?��e���ލ:i̟Qż����e���<���{�����/ԙk� !����`y������#��e)�������ҷX�5NSc�[�V4��I��	�Ƽ�Q�SQ[��ب����1?�ڟ�ڲRa�2��
�f�@�k`��V	���1+f�Xy�g�j�#^���TUm����d�-\�puå�[
����\c�\���w��7s��_a�wjG�v�~�����,CcaC~�w�^
�ѡ!��X?�j�_�ka�R,09ѩ?(����b>�p���X>�Q�a�hH�Ym@6��0�lpM��&����U�����\��p�����N��o`���!#3��:�w64�r�;SR�>srR��3K�I#x�P��B���A��(Udp���>��φ5�=����`+��J?���Pq55�	�k�ʔ������̙�M�>��˕��طv�R��֗�Q
 ~���Yh��F3�&{����E�u�?�U�m�[39�l%�zk���'��=����	�5�3�
�Z�� 3{IeC��]�<�|��ؠ���OQk�M)�#�[��)�D�θž�Wɇ:_hy����=�@�c���N?�M����р��s&�g�_5���	�?��3�A���{�<\�߀*���W����_�E#R����l
sE\��&��8�'.���o%������:����H��H���К�1g�XC�U_8��_����&�*M�