D�-6v�`B⧉����|j�s'H�Q����N��5�� +!y(������M:������Sk�֡�������).w�Pn�v���pH��$��Ԅ��hB `:� `u���<��W:�U?�n9�.�x8�d@c����.@����9��U�i9o�]w�����~�n6�̣��0���Z^a�^ٍ4�l5S�\R.�/�z��Pa+֒�\�#a4�9|� �A��p�;m��7�gN���,�j�Y>V�m�/���k�[J�`l������Êr��`�g�[�Sw�
�U��5�"�rr2U�jn�$W:��	�r2����U�fd(y!�0}�)�AGNd-	Q����/N����H���n�av[n �b�����9e�:_kN����ި��)��[�$f3?*�>�D��ſ*�@X���0�t��2�Ta�J��+G;�n��x�B�9v༘]a�|ı*�t�3�;,��:�����1�f���a�
�]�wg�T�����Ne����	��ڙf����̪��n�D�p7;�h��]���+Q_h�R����@��E�%%)JS������ə%aB��۽�,�s�v��,�Q�c��x-��|��{e���ߙ����s��{'x
���]F�k�@[}�TdP[���ӬJW܇r��EF���yU��
W�_0�r�\W��45S$@̕�d��b��qE�]KjU�U%�2��\n��X�T�����NVk�ʓ�0�݂T�ó�\��nxI��'��C�K-������(D�Գ��y��tzb:�WE�~j ����g�^;B��]��&�r-M��&�6�^���.6仿�$��0 �5�m/�,��p?�mD ʊ�U7�Y�X��^C39P7�]�B������	\�c��x�Pֆ���&j�2Cq�N�%^��A~t�����<��ne�	��mb8U0���D��\�H�^���E�\'�~y�X�t�A���U�HU1�ݬ�$_�q=ă����/wx��I2�����L�Nx"������R��en���� (Ke~��e��Yt�C++��o�\�9�v�x��������TdgϤt��ya�-x���ۏ�T`��l���S39�ϗ���T�������
����Y���L�Kb��*4�NT뒛�M�ð*>�=ix|���&�W��`����!��/��Yܻ������ҩS��~�)f��vQ�������of�]���=�����V|+yח���zݍ/f!8Q�R-�'�h؁4ZP@.Ǭ�
Øt��
H`:�,2�	����6���CL��O�?�f��qgeI!��e��uY��u5���T�� �� ��k�'�� �e8���i��P���.�3���@�Z`�vk�6���
qة\uO��v�a��E(�cL��!��?Sޙ��_aKj1�8�T�g��g��|A����#�j̒��Jrg笨�H�\f^N&��C4KM�9�U�|ԲuSU5c��,_'~�$sM��4���͒t�$3K�O�C�44Y!4ڎ�W��"�J뛘��Q�zC8ް�'!jO٨�~��+����Q�$�E�D����Q�7M��`�D"��^�%��$���|-�cb����ٕ�Xb�wv�m�!��m�G9��6-v	���C.x�rF�F�/C�1b�1Ur��f���8-Xߛ��@<���ry(�H;�5<�Ο9s%��� �+Q�}
��J�@��ʲ9�������%�+u�yu�j\�蔱��4�_;|��:�h&�;:E�6��ޞ�X4�:������oLm7΢�D1��8�f�`d��u'dE���y��<[�&;��t᭐��+R(��ȍ�d6�K���u�P G�1�����9`�dExV�mfvG���jG|�L��p9^�X.U@��K�5b��$����_�ދ�Q�|b��*J��A֐�lQv����h_d}r��O�*࿦l�xO���^��~��~U��W�Mr�5ϦdTN�qA��W���Ly����US�.]y�lP߁�WU|��7��L�R ��0ߵ�\sy1��eN�"���@��#�w&j��Ǿ���ٯ����U ̻?m�h�)����w�1����eM��{)g]���T��ֈs���v�1yD��E�8J`�p^y�F�F��,�	f�ت�8��>r��jR[^A���s�Q�����	-�Xl����y�������5%(b�J�ͧ������b��i|Y`p���zWо4Q�<�.�*�pK2���t��p���S���\��Q�
�#��Ʃ�yI]���Ux���r�8 
��Y��ݚ����;��32d8ne����*>�Z��X�Ǧ���49M�Tŝ>C�V�f��*j����ǩȠ�V�������twj���y�@����[<�a��ݝ�|�i>�c�^l����|F/0��<N�^SAup1�f��l���0_��#+��uZ�=���y�d�vP7f���o�1~ f�`����e����9ym�GsP6�'��G!!O��!����m6���g�h��*&�]TW�.����g�ܲ`�$��i�G�`<�%�]�k�ভK�ĝ��o���E�g���ۼ�hh�����w�2 �n]�Ncȣ	\y2@,N���%,���I2�5(�/d����΢!Ѐ�]׮1����DZ�^O��@��*X "�\��s|r�{�	���w�3�����s���:+~��_���ݭ�t!d��3�p���j���'���50\�
��YCW��>����-����=W2���7�;V�.�H��!�CXJ��������Os����s6���F�
	Z�˹�XQ*E�'n3��ɼ���QhX�)ǪZ��hh�L���.���!ۮv=<� �sOR�������yg#+�7���e����P��pe
9��<��T��TL1�����1A�&�vj�&9`�R�0�~���'����7J?ʑ�����h'�ߡ@���o��슽�`@����ZW���+()u��\�E9",�6pm�|�����D;Y�> gǇ��d��'ϻu����@!��'ՙs��1����n�f � �	vc�S� @#ƕ����Ii]���[4Իvo6��^z��ѥ��z߾m�Ji�4T8?zpY�����b+^6
�6��?��p�*���M�k2��p�b�I[IqX� �����#O���ĉ�Zenɘ����Fi^��-���m���򇹌��ܦ��©]���z�#�"�ߔ��{��)-��s��G����������w3���Y8$uD�����m�L�i��	��Y`n�<3�,��@ �޼��I��r�n��棛ݼ!��n�i��	x�K~��B�:���;��q�2�ą�'���f�(~�y��pI=�Hs�=��\S�N ���+OqiC�$#�gm���^')
�}^a�3��H�F����/09��0�h��SǴp�c����x�9y�.�����r�z�(���!�mh)�:�rZ��<�u8\����J&H�I����'�"	m��hjk���5C�"�L]%�d���}��<�r���`���P�3��6:E�W_�\�Ԁ��i,�ޏr�b:

�b�TX2�Y�0�đ<�R�Cd�*���n�I��յ�1�B��u�����7��i�z�X�E��jJ�z�#2@@;c5�.+�$�$�	�0��Ǝa�u���6-�H2����?��^��|�j(6e�m�>Y� g�g8�2j/�O��.�7�a��g;����)�_��ҮjK ���w8V_H��a��[k��<M����he(�!�&��Է5zSg����P��0Ң"r ���/gC�C{80v�P:���-+яL���Hĥ�իZ|��?�Q�zEr�֘ԬkW�w�%��B�p6NX������a
Ľ�4�R������N���y���͡4�ͯ(����C��H���UM�J:yF�f�Z�wsx�4f��m����WO�J�{N}��o�V�O��yc,Y��ɔr��/'/ֽ�=#	'n�ܴ�$}Y���ǤjQ����)�=m&�PW�d