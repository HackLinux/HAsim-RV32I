��0Vj�D�3l���ɏtҍ$��|겝9��1R�҇�ӗ'�9F��?��@��f'�d`u�v G������-�������&�+�0t	�qal���i(�4v�$��z&��A�2�0`���L��Mb��ߞ0�-��;r2 (/��Hә'��AɌ�%�A����͘�2�Wr^����`X�N�'zi����MI�����~��~u5��c�"���yN^\�1\�N�Ӱ���'�0�o���% >n:d���'L���3eB�[O��,�'	T��9�,��,$��4F���(��-��g^J�0�l�E�\�s^�s}��;��k�+�A����u%Fkp�o��Zh��>�������)`��Al��k�%%��i�}����K���7'���� U%/�B��� V�9�MA�5��u"|IF~�B|�[�,Đzv�5�,�_뽞<�e�9(�E���@��L��R�p�1=�
�X���b���5n�v ���	�ǚ��r����� �L�՚��='� 3J�+�9�v�v����	::�R�e��)\�,9��xr� ����T�ě���e�.�U\��_����3{`dD�]�*�Q�x]?�)����o2�H��V|m���1����\�3�
���Q�a��El�w:�H�j,K����lK >{d`��A��!̏T�'����
�x�\/��_��f/�4�A�Q����6~*j�5����k0�Ѻ�|$�{�d�r�	����WaCpXQ���� �-N0�z�T�V��+��s��<��O�#�LPΩ5ŝ���%��_t���uD�����4b����Ι��w���H����`/��̗rH6��H0�V��C��e�}�=���3� A�p�'
A�0P��Fd�vB�q��T��cL��K��e^�6���Zq7�W_eb�]����C�S�O���03ݸT�g�ؿ��L�!�,��
x�ȅfZ�/v�9;��qJ��`ͭ��  G���V��#W�v���:������Y,��@?�D�볣C:2�����;���	�kV��fL �ټc���X��L>�Tx���F�h!���ב���ǈ����r�x4��62 ��mrȋ��F���2pgv�����}�B��ϲ� bM��{��F07���¯6bPov�ץ����]�֕y$ �� ��vq���U�C݀k��EV�~���Q�!�ܟ�h������!�0|,��M�{87�6+��Q�W�v���5��|�Q�!�>V�?o�G�;���Q}j�jU�qw����ﱘ�{ �n��=d��tR�}nr�W�H�L��ށh�{rconC�?k����5�4dr��c��~���Z��=�)�ֈp�X4��L.*7��^���il��_�9s���*� L�# r�C���� R�h�oNv�m��C]O2b�m��~�,<(ѻ {sF��'z�~�@�,�$��5zYC�o|0rㄨ�W�;�u�d={oݺ������!�D�!"?��7�T,i�!^�����+�S�<k">LO|��-uR��2){P���.dSa����e�P�7�d3eN���/0�	J���"��$����x�����7��.�"�֒�WҔ�TS5�d�퐉�n?���fg<t}�>d�����'��f�_�zZ�ak�(�e�T	^}�� i8.8/h�q�o�-��B������~{\�5�5Q~&�����O��7M�V���-�%�ԀOjы�����E�բ%�K�c���Ƿ*��T�o
7�l�%����`�sW��`D4�k��K5�v���#�;�(���&hP�?�Dw����.�:)Wq���y5;ՂDI�sR�3��eDM��S��I�a�A�Q쒟.R�M����?�<�3��p��_��p��'C��:i��M�w/)U�#�X��0,����¡�b��ǲcP��}Μτ�L/(��;*2Nd	�o+s�+�kK(���w���d[����!���P�Lp�Q�1�7�v8|5����
�Vdy "�T/��NP;lu�ŧid��)��U�>��%���W&>)-�	�j��8���_�|��͏El`o&��y/���Y{�7^BP�m�,y�-�j[�����p�V�m�S������ݘ��k՘�����-�z2V�\z]?��Y��n���h��ׇ��Ɯ4Wù�7�ةkM����>lȿЈ�-�W��M�7~�����l\�S�5K��:�3�s|-�'u{q�Z`j!q�����Q��9�>������0|k�]�0oz��v2a|�t���V�+/��JUD�়�<˅

���_`���+ߘ���1�nz�Z�1��$~����9�O;B�6�q�<Nt��9'P�z�:��xr讒�S3į0�`��i\K({J���C!ܾ��T�޳:*���n����jl������T�Ż�_��i9��ij���0Փ�o��?�Uk��kz�!!�~ӥÒ��`���&;l�A	�w6�C�''�;��΄i+��xE[K2y��@w�����i�<֧{Vu�;�)w0p&s�F�(�b:�n�B�`�����x`���RƦl1���0�Fԛ��-�ac��	�;d݌�SV����z��l ��5o�a:�b��E����0́?�a��SI��f%�HN����;�o�`x�Hd��l�X��]~/��Yk(]�C�TΈX��M��7.�敋Ώ�١,_g|��	H6@�i7�m��ځyA�I6~j��t����BE .�䔽� xCjm|��o�>vNȨ����p:#]����B��������6��?gCX�xF�7���S�������k�8�9��r��g/������?�e!�˯-?�I�zbɌvv�h�D��A�	���e�,mX��-�4�Z����>ZOg�ZMb�ĥq������kli�M�|���0��8�,��6I9C�jB��4-�{��t�VjۖV+#�XT��g�ڗA���5k��R����ف�|h��lX�lX�m*&r���nV�&g+�Rx��ZYh\!�E���wc�Q��Wqނ���p�o#e���LmX���#�Y��@s���������Mm7���"��C��E�M�D�w�*5�������e?�y��v�P�#��t�#n�8��@�s����	�yeF�8�G���/���DW