�3PW����،�����?����W�~�a�_��     #2`4  Z  �?�1����w�[�{U�^��������ٮ�O���]wmޱ]� `H 	�P I�X�*O��A�A�$ �B !��*2    7�ܹ��}�z���0I$��������%P�-��{x�JR�(�r�Rr
�TW�� �Pt9��@F�*
EP0!
F��z}Rٷ&�If  ��TUY޹����Z���L���I�jS'(�j "�@�66�X?������0�m�*F��X @h�������Z�q���l� 2W�#u���m�7�����M��l���m�e��8��G��*�Hg��,�4����� 8څP��BBh�Kw��ZD�H�+Q$�4�KX��m5���*}<�_�0(KgW���qa��n���n��"kp�7U�邡�Y*Wܭ��.La�y�F�E�+؜|*�U̲��F����֌,�53)i<aP�ar�2����W@��� ǁQ�l���Y�ǅ���v4=K��)N���60o���� �H0��6k� NV��:�Je�lbaE`_q�B{�8̐1w�C	����"��'v�Hܘ-Oâ76%��� Z�aC�#쒈�6���wa}Fe����-�颵���{a%���3��e5�^�k�m�+�V`��[p�~��59����)3�J~7��4w Z)#uԶT�0�kr$��p�MT��j�H0*Udŉ�>�ߦK}�蚵tת�e��M5�e<�ʛl��}n�Ȥ��B�}��I��74a	`͇�"��p6Ù4VT��� �h: L&� ���1�4���4#\ۑl[J���1���Qa+�a���1��(�*aĻ`�c0\�!���"T��ް�%�h�Y�G�3K�jr�Ľ�w�۱�b�9���EgY�N������]�Lg����ί3�r�≑�Ħ�&&��琙q��<`����Q�`K6���e~��]\}����� �̹��?<������2ݷ�pL�:�uu��ۂ%�E���l+eA�I���6����X�~�?�婹�b2B����D�2�r��3N`*^Z6!"��_qf�R��5�?U�IO��5�ذ<��5��"궠�����\��J-���FFHy��Y8��G�W�sX��[~���#q��r�h`�V��IѶ2�cfS�zK}�.p#�l�5w����Yۆ�Y)$-��D�@FK6��B��=��YLg������q�a��W�r����<A��I��g*�Cf�\d�al3�J?�D��g�	A%駲��r��HE$Pl|�F3�'��[]+^��0�4��c�͝��}��i����|9ܸ�,�Zs*U��ǧ>�G�S�ׂ1Rg_��r\��!$S.��a,i���C[��<D!B XxL��BҊ1��	x�j��8P�vq�G�[(���?@�8�Ĉ��;̎�H�Z:	yr؋A
�T�(��*�)+��G��3� �mN'T��S��Z�҂x�M`�^���x�B�χU@�,q�"m�^s*X�0���t(�2�Ì(�@�0k���k�hO���:b��f(�_�=�X�a�E��.Za�!� �N���n�)�Q@����v}���y�&�#�����e��+y�1���K��^Yj�"�^
ى�!:�_`c���X:b�
����&�j؄F��`�����ؖNĬ?��3ᴶ����
{4��P ��H�ŉG p���}�����УX���\?$��n��M'�-�4��6��bi�M'���Q� �OY��K���H��B	 j��-=!���
�{�F���q%;Ͳ��,}��E}����J*lLL��\�9��xgZ����!����"%z-yb��:8�{�tq�]�2vSP��#>���+R,:�� ����4�
�RFrys����D2F>b�|C�N[4SG�����x�Ǆ�no�5J�b�u`]� �-���'�7�6����}��AD"gY�čJu��� ��;�'|����Mx������D�mQ�*�p�P��-�����P8�MZ&�4�X03����,�;)=�j�?y��N-�`�M�&jl��9�-�(�׳5h?H�4�9Ԉ���i�Vj�5���(HO�Ó�l��i�$�� -T�ŵ�5\�V�LN�!�ܡ�R�2(�vg�
vuo�8����8��2�#��9�20������.���-�\l����#�ET��0���OnɆ�C�O>�d�D��F���7�U��Sէ�	�;�#�8r�8�P�x=�XT7�Fp��VTa	zQ�� �GȪ�=�b�Y$I*�J��@�?�#��Q6֔^H,�2.�>b���z}m:�^:5>
R�"ȏTMl�N.\�� �xD�EǊ���������ڂ�����1��pB��/�Q&n�Z 0 �4�B��&`4%z�:C���N�Pe:�%I�Z0a�㬖EV��M՗~�c�L�c����aw ��1�D"���f.�O؜l��ua�)�NM"�0�T��)E��pxxqo��ol]%M�A$��F��_ªum{�n�*C0��e���v�1�uH���f4"&L���4��~q�ob��;`�@��H%�J���cffeJ��T�O�(�p��xlw�L;kÎ��Q8�p����������h�- �O1�s���š�f�h}[�Ζ�P�?�� �9�I�l���i/�n�n-��X�&�`�bT[��Z�n�S���,L����]�[~��r����͊��gr\�	�=�
9�)�%�|�"��@��^�)G�C��m��I#��k�
�7�57u�ҙ(�����<95�� ��|+3��`��d��XFN�W�[]�:i���Ld��grwy�-��QS�N�)p�Ĭ�9Z��\�4��r�R���m��8�+�m#E�)>�V���ub�����ԨTy��N��J+(�Q��I�`gh4�|J	H�ߖ��5n��|Y&~��tm�V�g��>6��NY��7G%ar�à��d҇.�C��ca�Ke"��(>#��������bQ�g^IP<y����c�sF�V���O�:q�+��8	F�;�y�*�!0�Gq:�5JV�,��:�5�/�O�f�KSYKz6��|mC-���Knh��N�v�����e�>��������1�3T}/�){��cV�l2W�h����/�]��E�(7�}v���Q���)Uwa?��䛆m�Ĳ� K�Ԣ��7+D�`$k*�����y�3C]���`J��_I2U����w��:]R�MDق<�fF�$DI�6\"a#�m����n\չ�rZ�6����x>kT�3gȧ��#"bcJH}�Y2>_`�F͈Α�`)2:HE2k*���M����%��]�H��3S0��u��lq�����Z�9��Vo�M���5=@g6�����Q#6��_���62��F���K}h8�τ�_m��+�{.�j�m��+Ϫ�,�yKPM:{�u�S0W+.���>>��hphg[K��~��H��m%�]j�1������Р�l��4�5��y��.}ȁ1�͟Q��iy�JY��YR��ՐO�Pѣ��X����j����GM㲼��>�nCY�oLgS�-<$�(V;8���!�����b��#A&�}6З�J.�9��]M.B܆�H�/�xD#�K2�b��9�k�b��8*�ʋ��A�����a{����K��Dܢ�v�E���"ϵe~���⚥ݬQhX�w^{�װ���HK��z����R�~<5�C�	�{�H\Jx��*��������k �{u��=$(��Z(Y�;��L�|X<;��v}Vц�:�6�z��z�w2z�(?ewEX���C8�������=�9!���5&gx���0B!�c�?/<*��3u�mKm���-�R�!=6��EMm<��(<$�x�IDdđ��4��wR�11Cb��y���V�D ��mI��j�\�䩋Qlm9��8��������ٞ��<,�7 c�!����&��&�l5�<M�+}�k$G�T��0�U�����/]ًN��Mm��\D�kx���~`~�]<.T_����Be̥TF�qP����%���,0���~P����J�k��Mbؘ<<�E.��M��R "�V"�ȃ:���'Q6\�q�:����O�������k�G�t��ϗ�ͯ�c 	��!5uK⋜�x���eS���󏒑Q���~���薜���@ ���M��*���q����+5Hy���ľ�os���8�j�מu��Gڵs�G!MF�ēـ���jc�E��<T�i�W���c�j�*?�g�b��7����dw��e��n�ju4�и��O�.���U6�n�7�L�����:�?�bd;P�)��r���~R5ʅ�>�`QR�1�-�׍T�����/eh:E
{��6/2%d��9�}b�N@�ᎩC7�(hH�|Q���(�������2�Ы�G�yz���D~	T�W�4Il��k0���Z	�����O�#�]eu:�<���9򄏳�(�~3r-���y<�hq<ݴG�2�7�U��,��2Hy؛1�ѥ0��!2`E���Vx�J!��t�Ə�(mUޙе�#٭m�Gݪ9ir���4��Ga���M�+>�� �(�5Bt&���>����Y�wҁ1���b�,�:ގy��ÓɓP٠�� 19����t2˷D��P�����ځBV�	��vP�"\�r��K��9�M_�e��<�J��~��P�҇$L�@�W
����%��J�a<y.���A#�P�ĥ�B�y��ԕu�t}�tig�����w2�p�H�����'�ƶ-�Jg�zV4*v�3�µ�c0��x�;6�z����՚/=�X#��r��W�$.4�é��8p��[2\U�[�n�t;��S�n��/c6��z��4���4��Vl���(��<h��[���z����ZnueS��~`m<$d�K�b�����ud�ֻVE��/gz�fƯgC�Td��A7���3(e2��d�F��Ó����Kx �k��_�谓9��f\�@�[���g��=����X}�Z�Z��S�����6K�h������������.qd9mT��N*x���,م����?�~�ne�~��v ��e�d�	؅�`^��I𦘬�Ml�)�'o$=? ]�ex��<f^ܷ��fX�݀��#��:[&���%����_�F�w�x�wlL�����,�s�p�}�`]��L���bA<���b0�D���4�[�W�^*�'��ʬQ���LIÔ̷��t�ыE��J82���bq���6�*8���5�[`T��<�B��b���l͜&�W7
�s���Y�?^T�=v^ҩ8*SQDBk�;(x!ϒ�$ha�0��ɸmt�UX{Á��������R���"������q�]�h�Kr��ZP��;����WьI��Ad�mu�>���Ҏ̊��yV�'c��wJj�m��C졐=�b��M�PdBO�t�L����89'Rs}����)��я��]T0�kB
>�!+h"��MG��G��D�+ 
���Q�3����3�yո̰|�o���Աz��El.�eg�ٕ_��0��$�J@��dP�}��J� �@���r��[`�	gi��]ώ���B��%�#����K�I�S^RH�W� ���Xt�;3����InI������S�U��^@�b��M�*������$?!!�"l��̪��&�VI���
,��������o�/Id�e_�����D�۩]�^�j!�&����s����)�_��i��8�=�E��N2�W�t��~��%]_�?F,���z�b�w���T���b�"d��wy�T��wy�=��P����p�����I�|���?�T�8?��Dn�<��*�#43�RpmP������9�N��y��x�)j�7}����VZB� �\۝vQ�B ��P����9@����e2���t|e�JM�ղo%s���<>��":�(�)Ydg���Ht��Q���L7��m"s���,��5g��-�\P��~��r�����̓6�ĈR��7�	j��ٴ�uo�O�:Hͭ��X�,ґ��\�
��5�G>9U]�v%������Q��VQ��_/g��h$��&N��N�3J|��Ǧ෕zK?��H	L��nW�$��◵���Ձ�V�೺�����;Ee�����>i�=b�na?��L]1���S;iHkʻ����Og�u!L���Pg�π?�'7"c#�CAf���oc�L5�������i���}phQ۵�;O�����0�A��i�"�*o���ԫQ�n��D��j��77��Xԡ���id7��Li�*��!��n+��B�i1�� � ��.G�gX�G R�8�pĤ�]Yا�o��K��tɯ���!��6�s##ɫ��J` �u�u�"��G�$�Eh~2m���1~c����,�A!eK�{#��C�PJ��P�!%��4)C�$8�0��Cm��ӆZ6B�]�@��gDk}'6�\Ȧxn��ץ�>��$��s���2�,Ҧ6�C��O�D}���WT��u�������Y�k���1��5iS��"sQ����&�<6���m ���b��S�R�P[��t��FLX|�$4�S�'g&8+1�JD�H��{� }��j9�ڭ�̙i
���8He٪�Bh$�+�(������XU�v�K~�����?by�c�G	�*wR��O��~(4���p���ng��+�+("�[�ii�}9�ZZ�aT۽��V�Wb��[p�Eh��M��R�	%�p�@W�4��CJ�u�u�m#^�g���W���f��w�mL�+�&��,�	��%f���ȩj� C~W���~p�cS���֤�<��5��d���y�5�Ԛ�dQ�+�;���W�r���0���# ���!�R�G�,����B?�e�R���Y�7T��(�\]�$����\yX���W��M��aH�n�i���"��ć�G@���>D�U��Ӛ{�JcC��é��(U� Q3ב�$�[B�2z�`#��2N�}mx��1���dr�r��"o�\ٞ+T�M��G.�-YVqXS�t����jO �b%D��I(}g�5��OVCH���P�HgέB[��CB�B���A#gC����b��6x��_�*�q!����$��@��x�D-���9���-�]Za�7]e�@�(�δg)ZhEY������^��L�[i����U�g�<�0n`�w	Q(c�1�b�l��j��;�}�CG]��ϵ�lG(��"p��%P�}�y�[1��DkrSr���Q���䵬�D&��$T��h��jϏ����aP�Ų�����4J����I��>��{��e%�ԁ�F5}S���B�z⻼D�q��+�+�@��s��O0�1� Ƶ�@f8�r���}W����á�*��Fn06����R,�xMD�����-H\����7�_�}GײֵM[#��@�C\�w���lN;�AiH��o��G��Vi��ƝG�'�L[�{���2�/E<B��Ó%���+k^�T�q]�v�}!G�,B���׊^�B�ip���y��7:l��l,�9+x�h�C@S�(Uy�a��M~}k�O�zY(���ZZ��^�8
["��`s,��B�;���K����^���5j��XO	5�k*�B�Y��bL�9v��&칅��2��(��B�H�1�^=J41>(
$�����k�8�v���A�z{�/?8�;��������+�md8�V�wWS����v�t��(0q�8͛�:��_j�ӿIb�F�sFx�s�p�����������\#*Q���R-'s��9e�<_Ǡ[���%J�*m��.^IGAV��4���Jx�^����f^ȿ����Ǫ�gv#g����
�X�l�����F*D�E*i\�g��%�{Ѷ�,:w .��:-Z�G"�h-�k����6��oEJ��޸]G�%�A8ȩ�b�|fA�`��Ov$p$���=m��!�	�����k���>@������O���~L�Y}$g�+��������vЊۢ]��w>8������7 ��iUW���#D5/��E��K��Z'NWY?B7TE`٘��!m4Ĥ�U�9Zp$z���kl�q	������f��p��G����s�8�eb����6i������>��%�*x�������[8�Cs�2��5������^��SrLZ<�ޥ�q�\D�/觉3�"^���*�M &�z*�\�2�(�-xwa��i{�q��|f��Aj��8&�����Lړ�2��m(��b�7����x�Ly.&�q9�"f��ؚ:�-��6Bɝ������>s/�(PǡDSF�=�[�j��ȞxkS�Y�}� �삐�-�՗b/]�6�&��9�ο�i��-ْ5C�<J���ą�v%���eT8���E��j�3�E=��Gr����2��؀~h��,Ӂ�9D9�)G�(S>�u�)�}�A?�e�����ѢƇJ�u⾻��(����iX��Xh놖i˗��v��1J(O �4�47���8��L�=��T�W��7�9���u���'`85/���8Y�L�ñ��h�ܦ�1���Ѱ�ѻ�Fk��و�:M�����xK.`[�yY��m�,?�L7=�G#s�uǙ��zF�6[��N�˅�R��e�����)�Կ]�5O��2�8���[Z����WGh����y�"w^E�eV�3�4���𥇴�]h�؋E������������}�X�PsVsg�j�y�/F�{�ͻ��^t'�̎#���uP����f[![УFP��@���|5��0�9u���y*��� �|=�Q�.�س��HOq�&�1��?�粩�i�Ƚ����<�a�K�zX�6��gY��Y���B����If��L0�H��B"���O�ڂ�����X�<���!����xh �	�Yg�:�by�	{:Һ��ʬ~�@��~9i��� )Ce�΍u>� z��4/�%Z;,\I�ҕ�L���]���H�xt���(��J�^׬�z��#����C�04�&��Om�9�^�p15d�����u�=��M��h�m_ԷFλm���� ]��75�rZ�vll�GU�ag�}�V�MTIΨ$�g���f�1u瓌^�k!v� I��$cT�/��j-�|�q��@����
��,6we�E���J�M��$�}��M�E=/~�H�t�s.w>A崄x)RZq��̻�׳�ٻgƊ`B+�Pj��ty�D��h�c�hf	��[{��7��8�	�\:�żӧi�@i��Z�?�e�U�W����������*%f=1�$S�BXs)��ɇ�!+�d4��&<��#�U��N���P��gP��x�g��2�̉ă�q�iɟ�RZx�Z�d��A
��p�T+"�l�5p֊@hC��mW��7��FW	d"Ǝ�(0��B��;��R�V�]q�Ȑz�ѿ�x��<┆N(�����0�@ s���s�������-ϩn�;�_8���0� �CK ��8?���ו����Ό�eC�v�H�C30��י-���Wu5�F6����!Z����bWY�^e�}��{+ȇ��ո��e�|f�S��N��q!��I���!�&k��H���x�^
� ���Y�q �� �	 ���1{G�4M����G�=���cB�		���<�eڛm�v�*���
\1}8���xۺ�K�٭b5��������eש戫���9�k��~�����"���c�A��������l��hN��󸞆�P�:QA�Br=F���f���&[K"m�x���{�G�$�������]�zR��QI���g�H�u��U��r�#c�l��񰙡P�lQ�����N�Y�Q���V��4BN�x������>, ��H��C�4��|�4@�!dv��Z�Z��D�p?��f�ZT��RΡ*��&�P$͹�!�[l�T��"_����_(<^V�ʠ5
م
�6X����|_ǝ�*Aѐ�ZdMb��B��"X_�a9ے_,Sbwv�n}�M�'����*�'=I0��e��!L׺(�
}z.n~!ɲ`:�)��%m��q�ϔbfO�qO��G�P!��Y�U4|�l��6����uSt�>�=�bBʨg%!�<��&�!A��n�<"�3u<F�,��˚�V�(D��Mb�XD<)T�2�C�lQQU�d7@� ������N(�����Ut���q���B0C��'9�#;!�K´�~<�E��9��� �#��S���Q¯��έ [|�FV0{?�i�	ԇ�3~¤��VT>��
	W	�D�Y�US���$e�����)j/t�M�Ts�t�U��b��R����٧��IT?O_ ;���X-���}��du�r���]C�B���&7�N�M�K���]',���.�i�y/�Gm}*�K_�sL�&NIUYJ��;G`�T�&��[Z�*2���uH}�N�T��b�5&�������~;�Z��x�-��R���:�
�� ������\Ѳ�(����Y��z'P�f*��b�i���n1/D���¸_ʸ�`Y���fK$7���1�.ޢ��@�;�<@�L�Ф�6*t�'Zm��@L[pQe�W[�O��H�S��"��GU����r�T�L�c�@�횓"=�9]j����`E�?8X�dq@�sXK��7�3iD�����5�-9	�W0�a��[]�]��Ρf����q3���onxM�{ӐNw�&C)� �%tOW�;b=H��bd��?/�ɶ�H[��b�����T�;F���
�Uk����m*`q�,�y�U=8��%�yg�5�5�N8��6�Y������ٰ��.��^UKy�g�������ׯ�"��������Mǩ�I5�FPF�h���I]��-�3"Ѵn#ɻ ��33�	9��l��<I�**�8:���zx	�ʬ�D�J�Մ&;�6YC��9� ��K��_�o]-͜��C�d��e:A*��A���\�<E����~a�u,�� �Ţ���[2�C
$�)%]ӷ�Ɗ"\��2\ܑ$sn^ώ�b�s��<0K�'���^/�����$�pw�4ɦ��S���4���o��\hhr�� Y�[�V(-P8b�,��;�2��|!�����|ʭ7[ӂ���9��vh�|���K���g����(��'U��O�lG˂��l�����I�A�ઙ�P�B�\C6 ّ���D���_[���W� ��J5nL"� �.|��\6�8��J��ȭM ���u�:�<��/4B����&�R�zI� ���F����I��4��]Mt.�5ޫ�d4q�e�	�1�|ǵ�W�lm�ϗ�h�A��n.��+��:ʃ��4�
`��ڍD{���Q]���Xˢ�
�K����|�_�o7�ˤUbY2��شb���}����x��gΣY�ӛB��26�nE3]44�H�>h�t$]����O��	~�Uq=��"�ͥ���5}g>/��i�RR��W� 2�3FNӔP���W���p@۠�%H� h��f��a�I�8����D;o��t�I
�ܼ@e�4���r�]G1Gj��G��������O�x7�8!�<"y�_�:7R���0�"��2�̊h�&s���jڌ7�z�t]�=2���I��L5��qo������ �1p�p��#����Iny�������<��]�	`��y#�H��LWW�c��+��ݲ�T/�
�����h��6Z��j�ޟ�א�	]FJ�J={y��kuM�-e�{p���oB�qu)���l�u�>I��{��<?2��Z~Nr�k��.��O:�*�W�D{����:=�ֽ��;H��fn��M�*s���F�t̫�B}  !�}X'P�������Ć�s��x�X,U��ṨaA�	�@W�ĳ�3�M�N�'�F�RAN31l��¯'��	{� (-X�솅<|s�U7��#��EuL��Sb�Wӡi�څ�~}$�/�4�����I�|�N��Td&\�b8�s�c�B`)F�i��v,@jAoG��D)��Ƥ�~�岖�������Er��]ɠ�����XGQ�8�W,�����=^1�NW���iqΥЙ��Q9�&͖�� ���a'ԻU�t�Q3C%�뺓��vzXm`ϼ[54�<���q��������4�d�vI�#�@�pj=P`_�J0ղ8F!ȋ�>T�` 	��E�f���r3y�o#��ISy�D3OG=gQ����s��vf��;��M�>όu�v���g����9z���Z� �k��-(�,�$-�Kچ�2b\�x�x��b�v��'u�؊�n{���9D,ш�9��Ԑ˷�|��%�/O����d�C:��8��7wc�~(
}RA�Q�wɾ %W7������8)�&���pJ�Ȳr?h��89��	�����+��-�����0*	8���R5�X٨-�H���u����`,��*b�����?FZz!��K�oi�Q<x"�f��t�Me�&���WG�q�%�>�s���H�X�`=��ɵ�N4DF�����.+F�4z�8G��)�]��>�I�?��@�5u��J�"X�t��A�s��߂��@�At&+�q���Ȩ�ae��_���;�3��N~]�wXk[+lF�h�<�K�年�o�2 6�X�wZ�Ᵽ��b�'��8d��`���P����̰�vu��ζJ*��H3��*�w����FڭxnK���4�h����=Gu<��Z%�����Z�q��-�z��Z�PY��C�)����	��X��[Xq�ߘϔՖ�E�t-���bb���Γx�
�e�q��dMr�3׆�	Q�0%�8^�#����Dj�^�9����;�C�m�H�B�&�S��#�AX�IQ *��P�C9���dݻ4�܋D���Ӂ<�Se�����G?_.Klyj���`��"�O��V�u?��Qj�e�ɲ��L&��{'d�g���u�>]�3nC\�ռ����
�f�Pd��� �R(a5(Q�zA��������{}ᘌ=�li�<�L/:E5wG��#f�>��m�$D,�4��[����W>��5��q$����f���6jD�e��h�g-�5L�h��f�}�b6t����S����RZ���A&p�_@7�:mi���`����z��α�&�L��!KtQWWm��:��X�j�sH�$�;%L&� ���O q��Fr$Z����H�lq��ϩ��A��xָ��$T_��f�+��m�Ce#� �.���&��\�>�Ճ�g^�!�ʰU`�V'7ϫ��0����	j������n�(U��X��@��M���Ttet�TĶ3�n�#��%@�+���|.��b����� ����XT�O93��!�
Mc��Ql6.�	R�^�ǓAq�d�@1�K� ���
<�]&������)�X>��46����9��ǟ�壚$/�\M_b{�z������_\[YE�eB!��ɕN5����џRr��qt�V<;�3���}�qr�'�����bT��@��N�{Pí�Iao܄?ڢ'�@l�Y��8��� ���'�QNB��T%�Ħ���垗��H��KjI�5B��� K�żg��1�<G`%�W����HAq>�2fҐ�H��n�����<�4`�)�.����m+8�ꡰDA&�a��F���� �LO}m��T�Т�s��B��V�bᤇ $m��bf�6�=9�r.��\�>lɿ�p�p�Y��&G�����O	�l�����//AJd�#+�d4]��̾�Hx��z &�F�¨Ddmş*��~JDΡZ&Ǵ�D� �Q��s��F����./��9����WB���ዣ4���\�d��>yڗ/��f�>G�g�ݣAJ���N�^��6� ���V8bc�T�[�nd���S~4o�%��-�9HS��N�1��Iۯ���R�]{�ʕ�3bڥ��+���Q�b��(���}A��_�!�����x�	hqI�
���g����?Ŏ0<)/,1:Ģ&%R<$�:�x���.V����lV��i���#���3���U����r��bB�[��0#MZAO�k�@�Ӛ�t7khCH��SXL"�1�	����+������T���e���(y�"C��
��"b�����g �V@|\��dP���w_�[*��`9�"�Zz��ӫO�(�Pd(��X?NɃ�G�sc���]�ȚZ��CE�B�Q2)��Rb�	�����auʢn���T��Q�~��Η���Yg�R+�n��Ʃ���f�TD:.U���2���TI��"�c��մ �~�L�u1cpgR8����[�Q�p��q-l��St!tj�Z.'GCI�p����	�t<��9�މHLơ�Ht�iI�9�
і���X��Pv.Ms�`Y�F�����\���-�@\%���e�=�.����}�	,�qu���1��[`��,�ϛ��L�OзHՔ*�!�wrx��^\吖Vӊ��f8	�����vz�����O�n��YF`�Y��$���>� [�Q��7ߘ�F�ƙ�w���",��:�$"�s������`o����}i�� �]!���6#J"�z�睨��4�݊�n��c��T<;I)i�N�q,��,O��`%a��A ���e0�F3h@ҵƁ7���1�i���?����g��S*͹���!��Δ�k$�e�|�46D�&�¼?�B@��YXG�͊�5�d��@���ۃ=�C��f �;3&�w�_e�!���0��M`M����ӂB�oA5G�gL:X(���kI���&�*��
a
���)�����Sa(9�ؒH6�*Gn.F<���:�c"���*?#]�߫6�&��il
�q��d�����-�Djc���o�7"��)��Mm�)J�@;x��T\�ئ\�ES�s	�[˼�k<5p�9�cF��_�Pt?ֲ �st=W�a���S�@�QZ3��s�h�Hrf��#}�t8�Dq��p���y��T_���e4cR������c9�e�uOV#�"�s�``�:�]��ex�;	�z��{m�k��}���PGD�聽�r���y&N��r2(���Ke�]��BZxiH�}� D�ʅ��J�0�`e�����ٛ�)4��ATl*G��?���_	������E���r �W�G>��%_%��M��Q�HR]H��VF`���AH`�Lsx�<�3�58�E�AF��Q��5�ͱ�lQu�)�h��=OO��W�Wd �X$6"�dn�VB(c�'��e�ɴ0���?fz�!	H�,�)`AC��`�BR��[FF�@
�����N���̦���5��p�7k<�w�Ⱦ��{����j4L���r4��x���@H8��G�����\H0\����猲XE����`���}��~!PWu^��ɸ�� ք����6�
æT{Ĳ%ſ<�~{o�S�����_a��o-�"��O�*��fmk��~���;xb���i�^
�k��TM��r��Ac���J�l0��� z�;��I)=u��ݓ�;��@B-�L��g�z]�X_s5T�\�:�qD6�*�/P��_�O��VAr�d9U1�*jY�"XP�=��#GĆ&Fy�#n8�J@s$N@���({��1��.�v=���hn:'���v>]ꝡ�BoCP	��,Iu���6#��u�O]P�F ��9u���%�/��,~�J"�u<&((���(�-�D�ܢ��ȋ��W4jޢ������3���0�o�ܨ��]��/����+���Kޱ�](��`�L�,���. Ra�HZs���)�0Ż��,6�5�$�ЭPT�y��̓`�_NZ[�/kWfC��.0d,gs٣y�e�Q\d�-�{cN�fs�nҵ�~n���E����U�q�kb9������(J=j�L�����[= |KeB���K��N�K����l�]X�v�t\�[MH\��� ?X-(VZ %\L�!<��]�*)%&Mk��[t�ȸ��3�ˮ���ʾP{���4� ���E�±�Һ�:*ֆUm&�����
X[�ըY�FZ�"bLj��L�.V�Wל�ܥ1�ǌ�WS 1���us6fff歬�1�5�J8��*&]Ŏ��FF{<[�~S�3�Z��^]��ҙM�6��L�(������������#�r/G�.���OH��2j�b�(�6��������Mf4A?\��:r��*Ԁ�k�~ܵ���.(�/��U@C�n+�ov��W}�T��9U�9w����q��Q ��9pO����~�<��g}���½�� ����}�N���\p�_f��3��F8����ap�\`�xg�z�7���f����=�����G>����!��G��9�_s��y[���~/�
{��������t_��~�d��q�q�}�BoR���y8Cy�{�� ��⤻E����_2{���y�Ə:�!�c^���>�8�Zɔt���7��P�'�D"o~Lm,t<�j#򂁓 �s>�j�⟍5W0k��JM���`��
^n�,	W���9o{�tg<��gJ�������|���߾��le`�������\�7y�\/G�4`[x�y�b.q��dA|��×>q��8���޳o������X��ػ\��O<E�E�&����\F�ٛ���/#����a)�S���T���w�������^s�۳"�P@N��w���خQy�Y��7mC�@��ˁe�Ed�(z>�R��.~5����2*�L}m�h5��c�%��C����o/��re��PY�͂�V�I���^!�[�?�狡���
M�N���麷}̯����؞}�d�9� �V���������B�+���Xr<x�����sPr��Oۍm(�1�!yQDuW�![�"n�Hpൡo<��8䘴8㼆Uo�I6(&��Qa���dٙ�2w��	�aV��-�E��eR���#MP2�"��m�ޑ*�{줃�X�N���T_ �������c�#���H���6�6���x
�i��
��$[y{��o����Ο�l��m=�	G������Bʉ��� �YɮaV��Ϻ�̀�B8o��4���#����)[c@�'K�<d$�Tg���,�@!yߙn��gᬿߞ�*Xv���:3\ :��j|ε�*���X�8Id�Wkق<�$�@\�H �x<���z�:��#{�znj=n����M'�B����.;+�2n�\��'$�S����!z:�o��5�!��[���,��� �]	?45� �'��k|����5�� �z���.k��ϋۦ�-!�ݷ�S]~"L-�vR���Sw8�;�11$�/�z�޵ೀ����F��N��vs�ڒ��@%�v��.b����{Cj�5��S�Υ�Sz�`�΀|CO�"��Sb�����u�{��[�Jy���d�iq�2���6����hb�z�<����\��[̵Ux��8V��1̊�}�0P�w�n6�~�kl����,�c1��H�������,ض�U;=]�#�l@8�<}�frLE"kg�I�i�qnv�����̤��٨ލ�GB@"�sWeE�ДR:p���g�>l��PR<����;cPc�6���*� ajn\<f��S9����f��}�%��}��\�ݸ�X��ۊ��X�h+��<h���|�6e+��5cR�M']���vM��M;s3�v��7Mvu��F;��]�CUE���&J]w���H�kcW������La��+/)�4r���c�!�!�:�~��hb��Ěq.�=Xޥ����t���r"���W�򮈚�����p�|@Ѵ7G9��0���I�7��!��'�ܤ��/+{�]ݰn5k��1h��߹�N���21��߼̝p�R��L� �Xo�	�;$�Ŧ#��m� �p���=\�F\��z���¿�������JV(���K���q��C�Gb�*��N|�!�E(��Q�13$�����A3K+�ў��nz������l"L�v# bc�k���W��[��Ё1-�i�?�I��u��?����P�m(Q��Y�I*z{j�t�" �xr����I7�v�i��MJ��}��[���`��QH��sM��C�_�U�Ҧq�$���%�-.q_M��(�/��S�P�_Y�tI�n�6�J��LK��%�]⳽�PS#M{�߳f̌o|�*�3C�L���V�)�����us�f�l ȵ�cSi֡���
c+OS
.��}\^~7]D���}�����H+����OyZ4�b�4QL��c�u=�>����X���� {ƮnCj(�*�YAz��f$*qGF$��A��+y��![��0�P�[�O��)	Hvl��=+����~I�6,�]+!]ݺ�IK���NC'}�t���8�1�������K13![w�����vwU�J8#�t�T�F 7+I[e�X"�"��Uq��u~�-���l����9���1L�`6>tx����d��)??=��:>��`�%��z�o��ULkL,u�U��:�j���7阚�_ �n�̿ٙ�o?�V�}�.�";�[����Pĕ_�&eW������ƎT�9�j�b�]�ƸE�v�}�E�y���uU�f�m�w�3N~�,�W�k����[��͹F����	#\��kϷ���'����*��l�a�s�ӱF��z�ui��(� �L����fan�D79�.T�,��t�/F֢�x��3�$7Ǭ࢝�n�v�.���Z��#����YFk�*e��!�14�ҏ�p�He݊����/��^uj�7�T�-[t?�������Ю����7�-�V��M6t�t5��(�J��n���6��j͚C���2��cS�8�u�Q[��@g����%�#9����z�T�z�`�6RV���o���e�db�d@�'~��e<\)�cm&�{��5�����8��K�xQNIq��d�)��b��a��B:A7�ks-4��Sgth��5�L~���9HbC(�Cv�պ�m�>�x�#��$\��BW�P-����;عG��;d�Uh�q�*��Pz��oYOmC&�؁[�!�x���
:�!/��j��?!ak
��%G\E�w�& �����s�%��I�Mܒid��e�OYz�^d���<O��J:��ێ�\1Q���n3n����ˇ���y�u�q���a��R�j���q���M(������%�Yd�!�D>�/3�Gl_��	��gE����h<l�ʚU��i��م�+��X���_Bk�;$V�v�h�	���R��5����=�\6�D�� Έ�����seX�R���HXz�-YY������p��>f)ݨ�l�f�-oT��Ҽl�~���Y$�`!j�O��~�T�T
��qU���h0wt�IUU-�\��j]�7����.	����WU͈r��n:�����X�����Us<uL�O�J��D:�]�����`����.W�9���X���'��/�Kӧ/��P��.��Qg�4o�����Wd�~�^P+�2����n��� Up�ݥ��ͩ�4��N+_���(�W�t[���iP�u��Ю��j��=5�ة�?�Hy�_����zi�_{���������@����\Dzqwa������������a�\qq�Ųl_v�^]������\Dwq�s݀�����zc�ػs`h8����Q�woǱz���k��8�Ȼ�3��Pw�{���ܳA�l<��ܽ���Ww�z��Êi;�q�۰�}x��]w i�G��;�C��aB��.C�wd��	R2���aYu���Bs�I�/�X�GjI���ҷ�z��0L{$�����3»��� z�l�`�aw���`�h��_�%M؋ #}���k���a��[�	��p�p��� 	}��ZT��ޱХ��?���}���7T���`J��^��.}��x�;~m�L�>�����K\r?��G��i�C���2�{���]���|�=������0|y��g�S��Y/�l7����7���<��������l�u���GJy�G��/���p��]֛d�~�8
~e�W���?�X0-s�3-�|�7ok�Ҧ���������o59�V��#���?_��p�1z�[�#����T~�ȿ�P����O��%�[��|��6k��>�o8�|V�ߖ���>��7����U��C{��x�2v�~��[�?���-�%>�������Zൗ��|�˟��o����z�y�?�w>�}���3�o����o8���w�����_~��C��7��{�'���n��g�rt/<۠of~��#��]|��-s�p�^z��Ʀ����c;���z|�k�ݍ����N|fgSG�M�g�H�c?�y'gֳ~�'�>��/�	�k~�_r�%�G=S��wҗ�����w�����/[+���bQ�~���>����w�Bẙ��O*|�j�)TM��T�_��;ܝ9v۞��}l���{�s}��^r�V3����}��?�?�>,��0_�nsI6[��2����FG��q[�n���v������G��˪?�O������A�t�"߭�����3ߺ�X
��Gj�é�������3_���S��ou=�s=������wj��O�S��� �� ��c��<��7���ſrپ���}�������}���C����,ޡ{q�ܫ�X�B�ƞy�l�=�{mGf㧻6���^h���n�+�+�����O.6�x�V�̯z�]�y�_�w?v�ozh���7�_д���olWӦJw��z��"���?�>����	?��?�,\���a���/�C�8�Q��Nk��١��y��/�����ܛ������Jy��/~��.����{O��V���ő�w����}O�$�H�v�'_�a���u�>��|��w;��6��3�=�ᇥZLq���j�8�Q����/8�y�3���Nն��ߛ�����A�ni�����׌����YWOȤ���տk����-�+i�z`G�}ͥo��i/�������>+�7��_��Z?��g��Gj����%z���˭V�q��\~���y�'��W��{�%����p�>���?T!����2��������u�>q��q�A�����)i����.1^���jy_ɷ.x�W��*�廏G���ﯨxg\�3G=�n��������ZTv�O�.���'���'������\ա��mٳ\����1I��������f=��ӽҦ�ϗ{ҟ}{ɋ_'N���}�Z���,V5.ֽ��U.s/?�?�^�yR�%}�+��������l�}����?����K���S��ߕ�����^4����1��b^˧��ٿ���cr����*R�j�M5��{r/M}���Jx�Ϟ�����s�-S}�۶��>�q�ܾ�]���{�==�'�XO~�	G��'5}}y��S�����˵�o��jf���ۑ���G��~��Z��R����/���W�������:�ȳ@z���N��j+������'~zyW��Q[�Ǖz���O���n�n���/���#���5W�O�A���=�w˸	����zS�ڋ�~m���.�[�/�U��[���g��ܟ��<���S�7��GX�Q9+����{Z�>�����h�֪���z��<��fW�|ֽ����RZ�vJ1��菦�N��|!�����-�k�6�[m���'���6�_3�O{���ɦ�e�R��z��i��F?�҇��Z���{+�3���P�>��w��k����i畾m�]���o�����~�5�=�ߋ������y~�?������v�of�8��������q~��xO*��z��_9�Q�����T3<VI���G�[5���_s{�g����;��O��>�-n��թ����S����7�y3���]��5�M�;��M�7�����񂟜���v�����e�eߞ��Nm�
�������;��?z�UjmGgg�ލy���ï��������]����~���WO|�/��m�;���V�F��o�2,���ߗ��3���i�y�;N�ԧ
ߜ?�o=����8c�-���﫼\�o�d�݉�y㮝���B��?ݙW���������_u�?��N�O�	���X9~yׇ���诊|�W�ڦ��_��>�ړ��=ԭ�����_�ߊ )��5RNq�n'a��N�m�G�cW�����N�j�a��c��>�ƽ���<%CT̸�P3a����v��ǧXyF�k
ZU����O�[������V�L*6�:F �ƕF�L�U�J)2������X�ժ*Y���*���V�L���Z|If^��[?̗�:j�LE8H�3ooJF2��#�����aU�b ����ʝv�y��ud�
���_1��I�;���G�۱6`Q��8�-�'K;�0��T�fd�cم�~-6�a\֪��=$���\���V3T5Ϊ�5}ٛW���k0vuh&���<)luj䊵���j��
v�J3�B�Kd�&�5V6^$�10�U��jIe����g��A�և�HJ�P�kVv�!wW���h�������� 	�i<�3aSmg3�hlɽ�A������<��:��_�+l�T]�����VO��������w�M��;�=�ߢN�����C=H�t�qAw
�����S�/pTh�cds{�̙%x�0d�V�îcV5e���� 	#b	É_�l��}���^�u�(sXXF������T�Z�7��I����FV����6�{Ջ� �YLwBBAǣnn�_,>(�ԴΖ���`:��� K��}.��f��R�c�/���=NT��
UD���JI���c���r���D�`��e����^�V���h�E�J \�Ol�$���d:��b���V=���h'��qDx��2��p}��_h������q6��o�_ǡ��_H�*���%�aɹO����e����]c|�ɝAfG�f��c������j����`��'1B�ћ���p��QkCF6$����b���U��ެʼFA!K��ES�S_o�L#���b)�E�uqځ1̾�RH��O��oBr�)�F������;�;Ȱ�E	�@�~���H^C���?̉D� �y�P�g�ƴ|_����� � "C�&  Y �1������1�o�8���
0REy�R;��~�+_S_�!���ۻ��n��n�ъLS}��>��P��p8�a l�����#�  ��t�JO��,����f�>���,��7ٓ1n�K�Rj_j�h���w9m>P��ʽ�I�B8D��-/@-U���SB�
��8��ϒR8�X6I��=�?  �! +�~{��޷��n�vv��I�\If��mn[��$��3�� �b&0x@UD�8�@�q�@�yu�s��{����i�֖�U���B�YC\W!eJXP�QuC��\�Q!��I(���;:=͗9���VW� �����^�̚�*id]:���G���Fcw"5��toR�����.�N�I-�ܽ;���L��~�	���{�uQ�T[Q���H�~���<��,dw����?ER)Z���y��i��)��`�+@B��;b
$"c�r(H��.L���@�HF�yf<|��T�d���HC����j�"2�^����}�~C t)�='�=߉.;x��ittd�.��$��#)�v�T�4!ɣ�������S)�!A��QӰӡ=�5�)o���T�ۑ� ��Qݝ\z�z*EJ�Ƙ�	����n�E��L����ä>5�ך���|ELL宯�������j;��$]}Ү7 8$��E��EK��N阊i��oק��R�(L�Q2���x �y���1M�^�GS�CE�A��;� K�,�[0dΠs���Ba%�,㺬��W�'�������)�R)�P��jx����jsn���6_bѝ�Ⓔ��C�����C$�������+E9*�TkL�CG��ф&� D��vK,��]�D�@I�P����q���Ճ֚}��D�GV��������M-�E��}�I��(�2|f�[���|��;�-�	�lT�&[��2�}�K�TMCG���A%��e�&#�tT���Nm�NE�D�+oZ�d�Qs?u )k��zJ��W
��*���Z��2��W��a�t2��Jw+S��y�(�D�*�X��%6���T��W�b	��>��y�{�#�z�m�wt1�>��t/�x_�M�j��0��
�8��A]���|��t���L$M��z#�Z�14[.�)O���wE:���ф����[�3�M�����t��Y�	�L���!���UP�&*P^nN+xN�[W&Dr��$.2�R�?��Fw���h�y���)�p]"b�3ΐʇ�غ�q�`YSlT�d/�ĉ��E������\���ց�T�T!@�0+X�E�D
���������=Y;��؈)�e@��.B�����65��dO�q�{g�@�_!G�^X˼1O��Ueq� ��Iz��^��aox����S^��DGKi�w8�f��]��M*c�(�,T��;n�+�����<vh�ϿI�<�V��E ��9Ox���>K�8��vX����������l�M8����{(O7h%_F$2Q�q������݀t�ly�a�m��D��\�����3�1�S�Y�E��P������]��#�l*b4�i���	��$Ǯ��!�U��sˈ$$r��4��p�J��8�2��vg������Vt���i ���W�]���}���o��w���$r��{�Y���\ �t{xp~�	I	Q���Y�2� �%�ёG(�[Tg�'����%���3n�	J�/R�X*R=�\�$y���GOFI�K��t�G��wؙ��iU��A�N.��G�FO�x̴q���l3y�r�xZf�����A�C%v�BN �E|MPn&M��~h>��$M[R��$�;,s��zU��Q��Q�� �D9P-u��e��4��������P�a;*))xb¢�U�S^~�Z_��)�=!��=R��*d�6��I��L���/�nE�υ��AF�FH��V��X� �˱M^�'�-4DT��\�{��G�uC���ga�/���;���AxEDTq�t�į�n�1~ﭰ�_�2�0�1N�j��Eg��ř!�,�w�s�o鿜j��B�2��n�	pQ���w��y�ߤ�"&�4q�ɀEP]aٸ�&�J	ڌ2*I�Id��J;�r7��Fh��{R&�fQ<��yRd5�#""��M\�7Z�2����91��"��C���z�&����[����p�F��Rc��m{;��H4�٫�o�oPl$i�a���D��:p���F���=���u�h@�����WoP$�l�i��P����	vM_ڝsv�7�0v�C���v�K;����v�C���9r9��s� �zwȺn���G��xL�@u'i�A�:9����#9��B�r j�"��\]�W��
{}D3b���������1�L0�v��K���t�,��ܝ�9�r��9�u
�u ��u�B}�{PR��.1jЁ�t�#[����:~#𘾨��f���ryw��7�a���taL�;^���)����?22a|"h����ϧ�:׉����0٩�L��u�S8cn�J����nx�]NZ��t>�{���ؚ��.�a �����`�6��J����x�u�"�n���|�C���Sk;�iZ���})Α�����|�Z���{��ӥ����G{_+ѝ=W*�S7Y��|Ѕe�9A���U6uߝ�^l��]�Fd��(NZJ�p�'"��6b?/Т�l���w5�q�qRǖ���9�DI��_WZ]6{�ﮕ��7v�{Zw�ٵ�?N���u�US/�OYըTS�����Ŗ-��ޱ9Ջ�>�8ۆ�}a�h���.|f7�Y�[�	�9g!_7ޝ�p�.����d�듷�ݫ���+)ZF4��r�|ͫe(��ln!�6O��������R����Y e8�NA�kUS������ߢ=R:��<OVc�v�B��H	�i� H�!�$�!�S+�.�W����X!�\�i�L �E�Mn���k��2�]�мW�|̙�usc�v4���=BN��A�ʚ.a���zpPQ*�%�BE�����{OMBOFMPe�]Y}�a)��."I4f_Ā���A+�[T�`��4�@O����F5-��u=���3;;���z�N�����ݞ�"ƕR0S�:��j�F���	��#���ɔ]"�F��\	
� ��-?3Ъ� �L��I��[�����0��~LI���xL��O��!��xک����@�Vё��~�"��6��Nr!4������#�8��A�N�h���j9�>ؚ�KTW/Q�R��:��C2�R[�H�E�7I�JVb��}��1P��N�Ѱ���I�	t�Ӊ��R�L۵��2� ��-���%�]b�F�eJٛ�K̫����CBO�]���~��ߓVH��Wi�f�Y��N��!��Z���P����@�,��	0��� I��싈/��0)�NQt�����C�b��'Q�)��m��m�Z��7������aU��S����B�ֳLJ��9���]����z��P�a ����eS�dZ�f�^=��g�㈬5�}������E���R8��<V�ww�1��T�'��o+�w<M���J�
��ٔ z$h�[��ȴ�;K���0��?J�R(�@���nغ�U�nz!�ax[5$��;����� ���=`{솨C��5Bxùb�<���B$�rOG�� �)td)�od����þ��Ɇc �dy���j��ߧ�T�k}��M��<�m�.g��ӦɩQ]r�86
L�2Ƃ;'���O�o�	i^��=��ŧ"s���W3�bM�-T�Q��,uZ4�=��pR(R�xsxV�D�D�[AV�;-D��������;6�N�ZRJ�����
Q�S2�bp�M�:�2�V2�� ���(�Қ�:j�+����v�=��ۀ�6��9J��;/�B����6K���i��6�����@�����Wd �J�O<�=�i��-��V�����@��s��~��6�u�n[����p'�n}8Ls�:nN�5}wh�i����;.FZԖ}��_n�� ���Sl��z�۶�i���o��Þ����S<�Hx��|�\j����^wp���N���-�Z�f���]�+^��𧞩�x7��.X�i�1;W��i�V[�ulb�u���c�h�_ҭ�c5��7Kު6w�1����Xո��-H�n�\a���t�����]�^jf��܏��ݟ��v���\���������ֽ����Z�ˬ��©|Z�6��������G�f�s6m���U�~�+��*�%7z��]U-�k��j����! 9[1�����+��R�S��i�-���[,ۭ����L�񙶭I�N��N��-v?FL���!P�4��cw�<�Q��*.zsy���� �7[�wT��{G�~��~��wQ���j}��A�3hShG�����<�>3_
;t��R��xQ�	b�L���T
��h�n�ٿ��C�0�.�j����^x\�Gԩт*e`,"�'��X�l�/�[z����	�#����O(�#$Q'�Qw�6��w�����U~�)����v���;��̪�:�-A���I.�Ļ�)�Q��YDZ���M�@q��k{C�}��ʥ�І�xk]�����$6
�S����J,ǜ�vh�����93J���~^���~��ݡ�{X��Z�D�Oܒʺ��aUfm �d���`q0���mt�S��q*I����}<��"")0c����Y�����aL���
2�\f��a��� �O{ ^�!�+����e4wm�Ŷ��2 ��PT�G cGJ�[�kd]�G[��T�,����������R�oK�p>nuy~�x��3�^_��,��+��m���aH)o}Ps�`q��`)��_Tvdw��X�%Pt�-C�x(��"��,B�*�`�׭�I0� ���|�r%PB�`�c#���V��
2"�gT�i�~$��n��	N���e\
hH�X���"��C03��i�29!,+-<�`�z�I}$ ���8AH�y��f��u�ܢ�Q/Ϲ	G?�p�a2�6ѴS��=8Ww]�t����O(�E�?��ʴ7[y>��1�C P�F�O
��[e��O�ݽ��wW��7[P����|��Sy��C��2���w�m��_Uɥ�{���}A
�,�l�QcoK!��ϯ����?��:� WD�α�5h#)�3ێ]���W�-�Y|�_��:����вN��x���ι����^�^٣��ǜh���zz�~~8�/�TqMń�/����]������BW�/>��囡����9�П���F����^�Πw���ᇋ`��̹�~�*��(B���`���({�Ʉ�\S��Pa�
yS��o/t#��M�����.CT���z#w^ׁ��^E�im"j��^?t�&�z~0 T�h�$w��O�B�;:xg�t��d}06�
d�ds�濡oV�.�A���SD�)��0��/9��-Ȭ��17[V�*e怪R�Tju��jű7�?.��=�@9�ꄲp��}�q��	�?�pS�O��f���.�����{��'ݛI���׀<=��p��;�>��W��G�O�u�oc�7юrΝS�����ӰC�y�mLnV�3�����;���I������!���>X����ue�@I�݊��B�U7;nC<��n��ٿ�Y連��v|�|��X��ۡ]�;�m�����l�����y�n�������6���}��j�7����~�
�Op7Б��Nܸ4fd*�7� E�W��7c�=@�۸���5�ӓh'��=��}z�0k��w�<�4���\��i`P/��4�|�%IL��w���'�Z�Fn]���s���`�Z�psHC%4�*h�C.�a���pD��l2�خ��V�a5A�ڬ@�6�+�$�AS����w��^�C���"&RB����H��Tdx�7@<t���1�HT�4�\��gT�ᨊ��שir/�ݽ�6��v�WUy����c��aj��Ч-�q*�[�mm/���5�>BO!��Tܻ��s�S�̈́�C^!,5��M�Y����VN=�TA��K�e8��E����Z�sw-��l�3��|�m5Y�S�]Ө��"�J�ɪH�*e��y���EU�����k�1�e;�hA� ���8�ԧ� oc�u���!ڝOar'�[~\u����[ϟ��|�8���1��rr�=�\�ٯz�׾l^��]QU-�vyn?k[8p]7خ#5Gu�ٮbV�n�M����ު�UaA=k�R�����La�p|ٞo����,6ƾ�ŮCz����-C��[��0�SD�h|�/��C����^��cZ3u��S'鈹�I�騱aQ/��=��*����˘
ړ���q.��(�h�ư(?j�T��Tʽ�!X�҆O���΅�÷�x�zKf�s��Gm��ʊ����G����[⛙-�����2_&���1� J�F ���׀Er(�q�JL3��gUW�Ye���`�Ҭ�h�/JL� |NG��#�V�]m��2D	r�A�w�T9���Q3\����1�]VeÆY�u#����`�e��r��eУFg�MXY$^�4�VX�F�q�����C�ނ%09��nMl\�Κu#�x���ĭ�	[�+3��R^�#�w���{]_@;�by�%^mX��Sڬ0�[3 ��?�sS�'����,Zs�u�cm�m��A��zE�n5��J[W0dF���uA^Q�m�\����P��Lۤ����x]�m힜�t�f�05ykP�*l�F����|�(4�q���qF��r�zq���B�.M��������)�d��NyDBi��^ցcP��,��5����϶F�B���]��*����j�Z5^��`J<^e�/u���L�@!W�!&��U0J�Y<zm�kc��6|�Z^ϙw�i�6R(���+E�U7��\�!���H�����@˽V2)��7�3 6d�`�X5��K'�xj�=�2��d%��ҜUޔ�膵��Sѝ�P���%*��NK��1�[�� ���m��ww[�rCֿ�[y��C�,�u�v�Vo�sXB�8P%UX�V P���0�(8����)��r�-�6�T�ҥ
�4�(���D��跟ڕ���y�����)�����Ǫ����Rd�v(��z¶�	r{���#����pS�Λ8@"6��
�+��5��tj'ֺ���~�@!�*楼��]��(��9ز�^����I������$�<ÂG�y`���+�Z[ �<'��@.�Q�#�5>p��2�ek�5��9v�2ښ�4�����ruw���ҡϔ�Bh���b��IXf�'|�E��ޣ���� ��Y�W�F�xH�;��e�+%���-N����
����:����~0gI�l��t��顸�*�Ƹ"��������WcKԄ^�y: �v��XC
0�q�Nc����xL�����$
�ME����F����-J=(w�f^�̖2�YQ��u�,����8��k)����<̩K'�5��)#H�y�K�G��M���â�YaV;GI/#�|I�G-�2��ߗ�z�����-rQ2j���q��G��W�-�Yr�5U��bN�j�j��p~���V	'�5����;:VhQ_Qf����)�q#�Miϝ�����+��|�	H��c���o`3v��\��{m�1��Ƽk�S�Mq��w���UNSO��6��aѯ2Y
��ub�r9�a#�.n�#�</p[���~N�nXC>x]旀ZB����5X�K��uzӗ*��)��K���,�4��(�B���Ʋ6mH��V��(�rT|z|���H��T��+�U���5o��nĔ��	�&&ff�*����7���rBD}�2~F���tj~����^�!+4B��ϼ;1?�[gL�/-��2�	�������ƈ��%���̲�^!Zg�I��Z�F�z?�BKۄ5�H�щ�"�W@]`���f��-0��G�����}U�&����z:�̚����r��9)���,��Ǭ�gEk荜�8�6���7/w����t^լ��A�;�'G�cL8N�m٧�^;�z~{�h�/�`1�NFY�����A �ѱ�T��N�3���Mw����,RM���g|��5Ja�h-������v���5�����=-��k��8!���p�����cT��oe0�#�\d�d$��3-2�*
�Т�$������fFU!��wU��&)P�u�����a�f�y��s�$���gX� U�_J,��Z�L��c&��_��5B���&<�4e��]A��-�3�	= �|�C�E-9�%&�m��F�&ns9>�>�ү�����*�!t��%���`��{��m���^sNE��V�`�t9�A:HxB��Y�3�^z�z�
÷=����8�c�H�lZ�R����<
o�ߤ&�g�c��8�F?�_��~`�%?;�/��֐'P�e<]e\�a�7�C5]2��[`����"�3&=�`|G������<^�	�̍����_RB^�/	4��D#����b�,g.؝$݀.I�O�/HK�}�& n��bI��3��T˿tP��\���|��# ��p~;yiG4� 3����?
e��*?����K�ZI��g�D�J�=�giv��m��;\��ݿ�	J�X;������'K�/�B0m	������D�`"���i���2E��@N��f`0	�#�x܈hٟ�3��MF�oA	�1G��x��4��As,jQV���=J�::�E�zIԎn���8��c*@J���
���~r��V�`�o��}��������ao�Zk��,�?��3��x	W2�Ľ?�<�(��9�������,��,�_��k�a�
M���.TT�/M�l�dpw��l�Zc $*������X�D�gq b`����>�*�t��@}Q�ҦҨz�0}�0,�Yj���	-�f��ww����2|@+�Y�}%̬�|%B(vS��^�ػ�l3
�'�����8�d()���!��/f>.2@�W1�?6�����v�X�;��~�i�[ M�+h!GK�~��>�eY��a��g�Ӗ����A��D����#�?2��	-��M�;�ľ���y�r����/�%ox��b�:8�Oӆ1ݫ��%(���a��lt��J���5�����*�;�����	]܌vb�@ϱhP1����ȇ�a����`]���]�]@�)��x"PD;T��>A`4_�,�͂#l��XF�\d���We�����ᱲ�w���+��FA��(O׷�Q�':ەwʮ%�Yq	��:��D��11�tٰ���u^)h���cx�?6��j@=ϟ��~TU?{�c�R�u?i(�]�Y��n�����u��;�����L{
0�x��jX�L@���]f2	�O� �`�\��0]C���,g�_��&��,:OrN���/�����1��] ���|A�8ث�虿����n�!2�Ek�G��Y��Eo� �i��ԝ��݈����x'�	�;up\Tˤc\x�lc 㴧Ԏ�������$fj֫�׻&��6���PP{�qQn��+1�.Њ���F���(�k����>P!��I�~k�N��S�_�F������FagTǳ}}7��i�u����׀��S���`h�Qq��ǥ�5�؍���N�X!�fx����|�A�xo�"㵠#���x�&>3c^�<�L;~�,�ԝuU� ǂ8�`��E��qn
��K4;-���o��1�v��u���CF�L���|��)xi� ����⫸e�ܙ�Ɛ�$H�bZ1iw6z����[DN@�ql���Op�̊����A������ǰT~�J��}��_��qkb�b��-��u0��oW�.9>w�@g�hm�a�(��	o�c�JK\Tx6�K��E�m5���)�$ǢP�v��>�������!�'���)�#&?��.�AjX���I�n(�*=�&���D8l��=Ӽ�hUes�A\ܸS�x�}��re)��-p�5[�C��7�����<.+��z�(���`ӽ�u�x�G�fz���ޟ{b�@<yG}8����A���+Ѵ�~=B�&���U��X	��f��>F�<64�7��8�ɻ@Ҙdb��Ǒ�2bv)삼/m'���}tl��S9a�u���q^����fdi�4�H��]O�z�V��;��Q���4�V�Ş��G��������o�WJc�/e p{� ���\�����fi�&��i�.���s7�$ޟ�=��c[zƥ���|1��AD�=.�P�G�<���P��h��
�0�
� 	xjn��l����T��g��q��_;��q� 
�ЬU���q��/�+$���
X��H΃8��Vf�b��"z�-�m�'AH~��`���hQ�T�˞�W���|��eL���]zp���J�j�j�~ߖ�� M��a٦���&�Y@��wZ z�f�#��ř�|2� �K�������$	Iګ
0c���&��y6��3ܤo_ ��@͹7�ж��5���x�<+�8�K>-5�~>��m����'	e��)���<Hf� ʗ"#�?�9ߚ��h�����Q�[�'O������1�jaE�1��,� 5��X��<��8:�Ͱ�c�e�Y�`���c�s/t
+\�=s37VSrl�QC9�Lњ"��hh�mֈ+���4Q9[B����؃�">2�)5+GgHW�P��!59�F�Ԣ��;�X�+���{���6��"#���e�͟����i�ɝ�������У(:��y\��k�8�
�����.R�gG�1���D;6L�fo�"�0pPb��KC�[�&�]�I�w?��<��z������Zy]fR�<`!��=t�G�XeDĈČtd��n�	:�_���:���݉c�j[�����nS���3�q������7�#ơ�b\�o��3��.W�W�;ƒ�$�'(��Il��x�+��(��+��k?�&�˵l���4��M��{W8���8��e�%h�:�%���� H�ѝ�R>���X]�@H��E�g�I�s7n� ����1�&�oa�~�p""�t�����͜��m�<��i�>�@ń/��hJo��@b�dB��h|��y�GS�T�`�6��f\*a��S���`(OI�2����Bd�������HQP6���o��i�b��+q����:��G���I�ʸqz���05��֢k�pM�me�k��"�8Lc���8�Ch(��u#K	���>����Y;F;9�x�u3ڞ~����ʜV~(��=�����P�aY_CF���i�����,��#-�7za45k&Cu���b�Րp�XM���f��Y�nNuZj�N����=��Vƛ5����_�,��Zc���Ma�d*���IU�H~�N���\�If2c�5T�����ЦP�_�!�/O�OEZWZ����Q6�^�C��5"[$�,�$�sֿK��C������x���r�9��^�1E����-����a{�0����7uӧ�28�����"�x>�V��x!a˲4�k��7R��$кG��4�[��LћcL�Cy?�	��]���ZA�w���M9y�~�4ٯ6�j�!
������@�7��H	��k�+�m�7}� ,��C����_zS�c���`x�3@ �|�����}����kg���_2%�
z'���ߠ�Zk��1c�Hp�{=2��`~&�`LzNU{�s���S�Hh{��S��`��rjC��4�C5jJه��4����&�'�fѮ���/8�0�5,Lc����+lΐLWu��L�M���׼Q��,����GYP���y��6;*��&���L���4�� �Bښ3�e�����8��EFON������&��H/��=!���<�����.��n�>���]Rt5���(%F�h���M��j����Wb���k����w>^q��_��p���� K<�\{���f���p#�9;kG�f�#�xF?]�~֜\XҠU�E��F� W쫙B���%@�3�8~B���lc�؋^C�J.S�*_I�$A+�J`:�>��Ԝ[��+H������	�����a�&9���8�4L	�K�/�p��&�P"�Oo�"��QI�b@�sW���'��BA�B�I��qY'��/#�VC�D�=�:���Jq�I�4�Vg|���S��f�s���5���\p�N�{��h��q�53p�S��3�J�}:�O_�nP?'UK4���� �����-�Ͽ�]����i�����8A!�.���ڜ�K�w��t��ށUg���]�Q�Ѓ�����rO8�ބ��?hs8$�Pm�ht|PJ���!o3�Ц�6,�����}7H�{47��B�4�l���ʻ�p��-�ECk<�ͽХ�wI�����%���wrw.�tՅ��у������}���~�����E�{�|� ��#2 V  @�Ƚ�/�ﻮ�_�_MXW���I�6��^t�8�6�lϵ]_��K�M�IDBIM��
H0*�TD�D :�3�"��#�E�����3�ti��hm���Ρ��.��e�.Ҷ�������v�ir`��KuS������){�S�]�>�V8Ã3TDx�y�DD"~eEVTPPT =@�V�Y��ֳ�����a1B;�f� W.��!�����y�Ȼ���(L˩#��{�S����=��Y���=X�)�p���u�4�*�
��M#%��n�R���)��ģ�����t=���,��[�jo�Ňle[��i� ����o
D��<���6�Yъ�0!BK���,;Ԁ�W���$lt?,T�?:���02�4��\����N�s3S�=�]�O3<�@-}���ǴM�yd�k2Y�{�����c؁L{v/E/=;���x�y}�,��p��u��oe���bD^䊪e_�ws6����|����ò�%������)�����֎��^C�%h�܉�~Rp������<������I�I��3�JGf|%.8�&����L,~, L�����'o�i����A}VE�N�<k}�l�K䍱fc,90Ooz�"��FOѲ�<E�_��꼃����~[��g'�h]?�$1Z��՘�h�3��g;��b
�XSv^Zٞ�G��i�Yv{d��fɸ�������T�%�=|\�0�s���sC�Y��*X1n3�뎖zk��:�=��0qt{�b=BT�C���a�j�E��F�8&A�Ђ���h.]VM���@��
�_��%�R�(����3S++ImH���u�Z��L=2	��ҹK��9F832ߨ�ƙ���bHM�Ť��&)?]��_�Ǿ/g��@��ţ�|JC2+mPv]�_[⾫�����)'L��%��cG��0h�]r���˝Á����s��YRG����ڐiJ{1����An�l?v����ڃ�ɢK1����])�2���ļ�@'�l �� �H�Ax�1�[��-��C�Gn�ٲ�݅)7q��x�,oڗ���a(�A���`mX1i7�����"����dN�H;	;B4�sO���#ﾱv������{<X�-�0߳�<�Z@�J�fu8�RO�PܬYљ�ñ�ۘ�Z��V� .zIj?��1���%�������F���z=?O�#�;V,���I$WhKW;E9BY��͑�fۚE�[�4�����[���Y�9��]�G�C�&y�!5۞=�#�����~�.?Ic�x�} U�Z���
��C�@tKd����?r�/�h��;�D��G��,<9�vj��i�����1���j�T
C��n1�0k�2D�B�}��_U5L��TL����P [��s���q\�I���#�+�y/�f"I+BN4q���+6$���d�dm�:�+K燱��@�E�8�K�V5R�#V�̩�b�V����X��s�j�:�%�yװA�~���vcxp�~ܰjR����O�]���"�԰�T�����0e{����OxS���@��ֹ�F�k����L.:#��3ƙL{��ٵ>�F�<�����{h�վw.XEί
�m�kޤ7�o��6vX�倦��z��rU;������<�^�adu<�����m����4��pΚ����xq�h;�j�$aS�L�\���u�Y�	������i��_.[g�ȩ�i1 �~B���!5V�sLD����������g��,�������r`�y�\��`c�[���(ut�쁤�dXH�{Cȭ�ѝL ]MECh�TjY;��I,���6u��ּ���1�K�|ۨ5�'��7җ�*���@�?��~����6Tn=�і�$c;��`�i?���IG��2�`O�Ųw�4�����WFQ���k
�2���/+��Ͻ���^m�fі���]�1�`a�JiI��v2�W���&/�X3��o�ZD�-�)����3̘���Qe���pY�F�o���J�09�=F���zW¨� ��U)�l����p8̌vO��1u���C�Du`F%Tۤ� ������?��qK6�Tn�����+�N�y�P�-ӻvq>W�zh��@ ���.ͫ4Sq�����^��~٤'�W�����p�"Q��.�s�>}��Go6z���ګ`'%��8_$A�=� �7�x�b�7ȝ�D�/��I�"�F-��>�/mIӽ��n�#Vp�2�2�wו:G�E ��U��y�ٱ)�u�}\ IJ�!Ҩ��81���ɳ���3F�JmM<TCNP.��q���)� �L)���,���sA���a�z��k��l���QQ�����~ls�n�e�Z"�r&�Z*�ӕi�����(=F"a�|VE|��t��=C�,9z 8��o���J����� 2�uE�6�/�N����e�(�
]Ň��k�_������Q����{e>@O���-w��&f�Љ\;�WL���<�m.���j۶/�=c�8�]���R���E���	Z����U9�g�!����T���oH�	���޴jj�k��i��(���.%�ӌpQ�k���ة��GG|˸� 4L`ՍќS%"%��2U_NP��_IgZ�����G��T�E|YO �T��'�nL��]q�%�ߣ�A��VɁ`�5|�J0����L�����L��uψηdw�aK�ۈRw���i��`$1�/HV�Wpg9(:'�:�o�lF9�<CRA���w�adɼ���ƞ��h�'#�����T@�Fh�a��c�ʀ'��
nW��Vi����s�ψb�Y5�ஶ�v�>�^����no8v O����]�(��������ì�	<�#��f��i7R�Ԉ���� ��uq�!v���?䝄{����
����[]&�?Q��<M��A���}Ih�	�ča<�L��
�d��vN�����5�p��-@��B�mieah�ʑ�:#8�� f0�D�Z�ԇF!q=ap�Fd����ƒ�0�RD-�s�D��wX�L��� ]�~H-D������z���@<�ߨo&r�Y��&��&�pd��}Zi(d�5�7�T0~�->6(���ؤ�r\ �k�L��iǛ���L`=���LRpj�cn(�ct-�\k����!y�t�����D��4�����q���UC�;���Qc��ůɁ.;�;%�x�]<�ۯ�"((��FI����ʛ4���['8��-+j�8f+y�%����wî'��,~$�[�Z6ݩ�<_>qB�#��:@�	$�y��Z<穟=Q�ün�WLE��?�ב0�)���U(��|�UԨ]YĹw�VC�VX��{�b?�7��7)s,�A��	S������ZBG�x����|��i�*�@k~�diio��%m]6�q�sY��E	��=F����ν�l�Ŝ1�]�s�K�S%i�TvE�Gm�0���������`�I^:��+)b��W#�p�+���+g^�˔g��]�eh�DR��^a�O�ꭥO;�j\�'��*�h��n���q��@Ѽ�J������cA�]�Q�1�a��@�������r��@���ht��ŎbĆLe@���(��y�00Ր�Hќ��GT '|O����c.���T15�i�|�:�+�qXi���O��cg�6�]��s@Y~I�R�^�N� �i�y>���R��;cw�z�4�MR����E�;>O��銩�F ��=ţ~\�C)�� O@-�\O��.��r�ix���պR�}���W��zn�m8#��oV2�S�dC� !�=�#��O���B�x��[�E�_��A5�el��x�1G�^6�i�sd�ת�e�W�i��b٩�3HO�@����V��˳dNR�W��YW�|�0����*8���R�q��|�[uq��< ������ն_��/�橠qX'�"D<�����Ō�%��׋b��W��(NUX��{,쁒|a5ԃ���	�8��T�����$k�������#��S�n�=r�@s]u=����ʼ�F�J��~GG�/e�~Ͼ�ָ#͏�檪�1C��ұj,4�I%鋓2e�WΝ/�?8Y=R�r�҇]Y���>����O�ꄨ�׮}��k�uO���=�WWm��\��RlD��8э/�I�_��9���{��m�i@K�e��b��7֎b[萨7� mIpU��kz.���z=�Ym�]��-�i�LAn�؜�{m�z�u�j��I =�x��{\�Sk�O��F)4�x%}*��Q����A~�`�ޕ�ʝն"ef�P+*�H�}���s���܋�x�l+����zc�UQ�?f�@���5ˮO��{œ���*vv{���Qp�&�/�^��z��l�{y���e�W�Y�ɧ���5l(�_���W�IX��/���W���1�2;T������K<�����]a[��F����W�<K�8���)����{����y���L������ש�{���巟�'���݄a��������.�_������a��sw�����S���uI���߹,����l�>�y��{�Y����Tb�����YnmnY�o�1`��o�璿��ŀ��g#�#����v��t�r������A@��D����o��
���~�����7�u4��+�/�����'���?���o.���i��kk�O�g�߉� �        ? Jy�7x�B)W.!�(��.�/q�^B�K��x�0*"��R��P*���   �U�n�˲lme$��LmN3��I�$��E��"��|�=�(ڕ��G�Z�]��t-��A/t(E�ؘ^�����n�0�f^i-� �  3f6 �����=�o��|���ڳb�IŵձM�X.Eʀ+XE9l�C� B� ����#�<Gxx�y�y�����zr���z٨�I�kqb�pT�]���&+��MIDY�
o�+-.��'TT=�+���[�O�T6#M������L�ZFY^����?���wN#u(Fg3�@�@���	�J|��NJ
j<�����8�z_��Ap�|�WX��| k�Uzw�"�砿�+3#s�	�w�H���q̧�����MKQzРC	��g����БR����5�9��K�ڛ��4�<���V����'Fh)P
�j2�Ҋ�-sUG�iQp��Y����"���Z�5���% ��Do�y[��^�26�s�@W�[)�����.fz�BG��!���=%��G�D��֜%�p�}p���`�`z��k���߿w���~�kM��@��0˧,.��{k?~_\�����A{�A�����k��������֓Kwڔ��i$H=4|�K��T_m�r+؛I^�����şoK��1�qn�}7�*�,d��(�㥧g`{�v%���N����}���^�j��o�����~q�J<�w�=��7J9r�~�n�;����=ܿ�����Y�)������H�{��4���v�k�U��_7�3�$7�
������LzFw��F�%ZRPOe�5mu%Om����Ւ��N��IXIZ��j����u����,���!7�EP�������c�����w��@g���L����pӆ��WP�"�_��A�{�sf�^�s��_�d`�6�!��� y�W?q5=��_}�+�P�@H��]e��U�`�B_W�%>P<��v93r�_�6����4��|�7^���8	�~A�}���7�I�?ۀ�?�	V�Oi �N���;�����bx��ܣ��+�.��Z��(�{����9$���m�!��^�l��ws���'<�WQ8s������)!<��+ӏ>5����o_W�;�%��7�%mo��S���w�����54����~_��.,x�sg���v�~N�N.^S��~��5���$�'��B"X�	�!
`h0ߕyE+�F+�.��!����,�-��]}��}�o-��X6���yj��I�~��CdPo�����h�WV+����{�z��� �CK ��aDOY/�̕���e0���������~?m~m��&@���ȃi����� =��*������[y;���&������������|�75ߍMise�,c(U��D��L����[r�_�LO̽������ǹ��{�Ղ�[�N϶|���T����Q??��b
A��
\���[�Gt����;7����1��K��0���"��{�� ��?�.Nn�?g�/�}��<�k�3�)���hΚ�����/ī���"�g|P|_Iy�Wf#��3>��F�P�V���t�_`����'(>��i����2>�SU���r�R״��$�t�k�M�T��g�@߃�z��t
�S�������oFb��
�K_����f��/�^����VS�R�S�/���~�����z��w��sr2�(���&�UO��i8������@-./sxc�?3��}�C�Pz>�g��?�K��<����l���S�0��+��_g�6I���̹_�7K
�K��Wě���7��y�07�P�W��>�Cm�K������K�f���|��9���</o>9�WD�m��o}W9^2�l���oWu7m�v>;o�k�W{^��S�O��>��~��g����c�_��0�WW��n���W0����+��A,(ض	!�V��vp����6�{
:F�\�p�	t���qG�A<�!h硣)��h����m{륽|>5դS�ސ��Qx;g�Ѩ*P!G5s��(�XdM���/��q�˫�#��9��VgMq������Z"�풴|��n(���e|������t,�8S5�;#)t$�֒�'h?��*��Y�R�;@�Uh��r#(d�#�]"«��>�#Z�ǜP%8���ɲˑ�62;w$8��%�-}���G���m�(�`i3�����bL��"��rE^ّ`[k|F<��wRw8��5���#���$,�S����l�G[��X,�kn��&Z Ą#)P ��.�YYF3�&^�UVg]�Ӓ����C���h�C��2�z�
[��`4�PE��;�k�9b�
���^�ˬ�Z�H���J��]=qɊ�e��a�Ip� ~>C$4�2iM�i��7u)��<�q�����8���$PKn���U���)i�� �K�kBu���C��KH��V�G�W&�� m���:K��n���c� 'g��X~�)&WZ���4I�^� ��=�4������^F��/���L�o�2�3��h��RM_+t,�d^�9�g+�:ḫN�r�.@h�Ո��&�G͜�q~<�I@����S@���R�"�EV�I�Z&cb��	8�i&)�����=]��בE��!Z
֥���υ؆�sN�Y�Ω��P������M�t���>�>K���2�ƅ�\��@��$����\�̚�6���!���R{�V|� �r�6��<ݵ|���i��Zn)��Ύc��O�L
��ǰ2��[��^F(~-��
l�UW� �7��][4���gҺMh��-�ȕ�$�x�r.�H��e#1X�#X��S�Z�9�ׄ�����H�D{�k�p�
����a�Mr�*�3�^@EȀ@k^�V�����1��յ�O��bMA���p���z��~�>���x�0���0�ߪ�)@k]�Ӗ"Q���Т���[�2)�H�����gAÛI�!�+܁��c�Y�hd;�dvƞ(g2� w���7�8���sR�M-T�p�����s�L��N-r���6� $�[W��w-ҨMh���.K�b��V8��Ij�K�@)V b����b+��#|�.B�_j:Ⱦ&<�y��I�=ܥ$�Lm�Ox0a�pIo��j�&
n�sP5�sr�DZ�P�g��Bj�:�W���¹l��1p�o���)�_j��aߧTg[r�b�~t뢜Li�yE�N��rԭX2�r�]�����P�:K�F`.�i�"����;#���k�]��T_!n�r���Nx1P�bM�U4U/P++S�i��C�F����5�t�-e�lk�͎ �3�c��6�D�.���Q��㶌�/i0
딸E5�@�a�����9������um��s�\V[�m�6���O��46G�wy�E���ؚ�QߠvqWN�F�Y��$S'2T(�L��}\�*D�/3��� Ր�l)�Ú K�	�:�ʤ;٢����dS%=ɛ�7hN�\��T��6��[����=�W�O�A����@������ R2��k,ok��?��ev˙免i���8�q��s��a'�a�BQJ�m�F(�$�5�a��p)�D#q����kPĘb�"��[��/s��MF�8���摣�tdiCMp�7�Zȓ{L��M1A6d�PZ2�u@9��R�0�!O�m��'��`��ܡ	�2(k
��7�������R���gP1[���۹r�����z.�śӘ�F��ˬxÃ���@v�b�t�$��w����p�1x�u�,��ay�������{lO�@v����4�\5K�`�`UE��]dr�y�	"�Ԓn���5m��/JR�'��6ʹ��Ȓ��M�����TU�� K���T�<��t4C��},V%���v��T� �p�Io�Ѻ�g�; X����~��/X�~��`�`mh?��Ƞ��- ߄�]G�ۻӎ���0������!���v跎O[qy��OK��֨�Wx��'� >q��pbc���������Kuy0�I�d����5��d��x�6��(����m����,y[U�V����_��B�~U|/W|M�%Ԝ8���%�GB,#�dѶ�u��K�Y����L!��{:��({Ae����o���j���bY�����K�~:yd2��ɚ�I�ڵ��wPT7�A��>��{a6ߦNg\cW01�z�X��Q�=&���3�Ě����4z���M�\y}��)����%�`�m���:��������M�{&�q߼�UXrrߛ�H�"�������(��>����g!g����KggM1�h�ذ�Y4���ab�+. ���P����|da4_�^�4/,��+�k���}��~��������9h&a���U��L�-r��/"�ߙ^@}����F���6�)w�]j�[�q�6o�����!�=9�g�em��#rT��*#OO���*�O��Bz�͞"����g��Sa<����Rvb�¶��}����W9u/M9Đ�a�/��V�����]�=H���=���Q��%�M��a�~��_,����������a��W�CJA�Jef�}I�H��'��~/s5ϵ4��_>�{���
r����<�����Ʊ�;�<���N�;��ſ�6�CO����$�.�0�wt?��u|&��y~���G�"�+��~�<�P��[f�?�M}�RD�l��ka~���I���§,��?b�¹����.J��P��a��)%��[�~�_��i����=?�S�
W�	d���Ϝd#�0��?�>�0򸔣�j?�A|�GK?�'zU�;s(w	G�>�{9���Vu�1�Ď[@���w���U��_�Aϫ?���ow�:_af�+^�)����M��؇�֮��Z�n���g�z������x�JR�wb����3/<��=�����ꮞ��� j)��#c�+驎�G�k�s������߂OLU���d��{��͌�'i�8ڽݯR��?$�<e�7�}N_��_;�uO��ҁ��.������[��>�N�Au����X?A�E4������\Z@��y��o�L��G�I��gf���AT��>���Qo^S�P�|�+�����\��O��]�=�������5Ͼ"I��y9����m�\��<��ғN�����?]�(�Ի���[��K�j������c>N�y�g�{y*���;���s��h�����o��@�!{��XFT��ˊ�Q6�H�Y��W�J�صغ��ZyK&�WR(iN�����ﾢk+Mۆ3p�`�%�����u(�GR�a,=�l��CLwP��|7*s�������ִd�CN!ÛB�
k�~x�d-�da����}�v�Ug#�`堸������H�I�Hyͻ���5�T!;(ϩ\a���.&�[5��n}�cj�y����3�C��B�U�U,)�V�ī:yv�>��b�2��\�bKl�@{q��|��t�C�P���Ӛ)]`Y��8� ���ZZ�T�.�P@�q��oK��lΰW�#x�hص#5��&�l�r�@"b���t&&U��g�Ѱ"��U?(Kh��a�c;��
�j:�Ⱦ�_��p�h����gS�r Q)�D�©��j��p�H�xW�B��c�V�e�ԬÉ�����I
?a�m�f�)�ŵ�P(.Z0/~SiĆ�a�Vx�ZJ%���cOU��:=q8��W�Y�J�:7L6n���4��#�\��Q{T ��s��~���Jq<@�i�I�[�M��p�{��U��d���/��Z��Ѓ4ߟ��qHX�d�{t����1t����~��Y;�K�B��*�%�/E�j���QS�K��dn��:��<��(�b:DcGS~y
��],�龒�׌�A.�]���㨗9c����ղ����a1�g-Vw�i0Vm;���%�W{$�@��.�N�͵����GHdcB=�NB߁Q:y$3��("�ő��2LA��HK=�:,�P��g��(��I|�S*I�z�f(�+J��I�1�խ�9߁@ݒ�Mc=�3&��rW!\���V4G�S<��MS���]�s7�7���gz�\j�Ndl^ύtP��h���q97�T֮����x����d���L�9���&0�w�Yg�KM���O=*$Y��a��/�x�C��SA����dNq��-�"�N�@T�~<�!����w8S�,�Tk3n��7a��8'���~���zx)���F�rA9w��5eCc�5,EHY���#�#آ�}�v\�C�B$c�q� NZ�\x}�Xj�S`��L{ݐde�p��\� �;t{��5�(5Q�Ք��U`qý[;�Iƍr�Y����@ɫu�O�R�{�ZK�����	���D��EB=�͹훛�HT5(5��C18>f�3�Ӻ�V��M(����N������n-�N�b��q��i�����#��$>N��*�-���/y~�j$�*"~��@�cC�T�G�P�J�'��wA��R�qNw� �U�wӞe�E�q[�HMX�(-[A��x��Fc��!>�I[΅4Ț�3�J�l�1c([ࣤ�n7�3�93�p���v�R�#�kœ��l��j�������j�'a��a�,!�be��=��U���7v�G��J²ܘ�zD���ta'� ��yǭ����[�БHFH!��2�?�U�9��;�E�v�mF��M�R����6hYY;�A;h�����\N����m���9�#	H�����X���*����zԛ�c�ٌF)�����KX�ſ��ÇȈ( 1��0XZA{�|�e"�B팺d��ۓP���4��9j�M�|~555��{DqwK7���n��\�5'���M4�k�����t�,H(#��g�br;�Љ�M[h$*�L�Ϗ�����w�e'x�u"�T�;qko�Cx����Ѹ�`՝�/B �lhF���E����懩�M��#g�O��U:��Xu ���Ay ��J:9~�Bȉd�T:j�>`������6M��ȷAg��� d�}�A�n�F�墘[�-���h�ze���|u�>7Mfi5�=9��w�t������&,�nTQ(�WZ_���xI�4Q,���Ǿ�!ƫ?�D^o�������ԙ>��k�2��1�#[�g����^�<g�bp�Ng���p�x��k��Dh��΢6��9����5i�*b"�t��#��/��`�0\p��B7��S�|x�����K�	�DddND�n8�b��NK)����6 �mN��n��|3�gu's��v`�<�-K�ښ��aQ�d8�i"�V@��=G%#��a�9�uՆl�m�K��ַ ��@sm0 �ʬDNA�.�'����cx����܃��Nc �X<*hސwf>έ`�W��`p����}�I�NY�ƭn]#�ԯ\����[37��i�S܉n�	��y�~\;&W�,2���6��k�j3���'a�*��׬0��.󶩭x��ܹ.�=^���e, �C���7�����F#���٪� [�3
$��;U�`Y�,S�a-T��7�cR�+��C8��G5�b����Z̑`�zED�@�z�q�����pz��E�業�fs3�!�V�=o�jϒ}M�I�dU��b��}9N�"=;�l������� ��!d�@��2+,�Y��W��i�Ӓ�l9���ۃ��}�ti��R��]5��b�XP�t�aͭٙ�6������	xCC�(n�ـY�n:Z��������Ana� �^��(49@�
��뻘�h���Յ>��z��6���ޚBG�І/��g8X[%�̳S#,W�m2�I�LMG�Y��n�H��zk�M�� �[ڠ��|�y"�(d�8��J�Fl@��hG�2��\�K��sb�qmn:i2$�u���ͪ��ˀz�bZ�mM]n�ׅf+��DSв��$�h��{U��j?���N��r�21�&}&�8_r���5���&3�Z���ɕ�������C���F�D�j1�.`N��Ƅ��[��ɉ�Z.�C���ދ�H`�C��Djq����>�g/Fi-3?2.�ĳ�l�Z/w7�r�Q��F!r��Z@���&N�xP#�O �{Uv8>�je��]d)�v?��g`+Zs�1�t��婎G�G�X�dr�/X� ,?*�Z�c4N7��|��}I��!3�����F���u��ǹf��X	Fzp1�c�:�Q���k�
SP}g��<J�����#
�[S�[8�2\�������<$�Uh�#�ff�����i��M�͸�X��DQ�[��41�$G'�w��j�OVU�: ��-�.�>^��f�pÄ����!C2�Hu~z+�Ņ3�
	@�gn`�WI]����ނ[3KI�C%��oх��l@Q��z/z���q89Eb~;9����B�A��n����P4ao���ug[%�0W��6㱾*��%V;?ؼP`���0=L�]`b\^cab0Eb��~�+$����7l¡D�u��a/�b��U03Z�x8eH���`��=#�z���:<ce�F$R�82&L �KӋ�-z���� [-;���>��3�v*�.������n��sG;���D@������W�oJQæ�9R۟�A[��K5�����iK���C��Q�,�(J��M;��\��@$��u"x�C�,~�ֽ͢&���;�
7$b�!T�*�^G�իT���c�.�ѱ�m$7f�n7Z� ���q�8���rfx@1CZ�5���~y���B�>YW��A�W�g��q�D�bv��0І��^�jp��Y��[T��NiG
Y{�ب��F��q���#�e��E�S�6����%3.��|;h;J�|{�Aj�T��F���'��'TKj_�� I�l�o�@1r�11tsy\�L�gr��V �,���o��T�����i���k�������I�%䪴
G,ri9�iÌ,�:�C�zhY<kF4-�?2��.Y&Z�}#]/U�KF����4�y8����a��:��V/Lf�6�y"0;S�|�v3#�[ݗ%hd�w�9���f��5�ȅ`��'��s���������ܲ��H��|-���D\�S��a����'|{����J��O���A������|���}x��@����:�����r��܏;\`<�I����d࿡W�}�9����?��]�w��,A���.���z	��A���g��n^�?��#�`�~yy ��ӏ�T�:�SGTA;y�xXS#�#6���ޛ���G��sȝ��y=��zO�r韂����g��wr�����p�~��ޚT�?i5���!�¤��/�tM��=o%W��֟�4[6���:4S�?��aqn��{��������A���=�X�.����B4���w���^���~��;�]��L���1ܥ�Qs�`�{���������@9A��Z���,��=��]��+V��~Sx��7����3�����]�z��'�gÄ �u3�R�=�8�^�w���"��R;8����w��t��w�I�	����g���?����_�R�#C�#��׬���f/�N�1���
ݚ��������ӛ/�5G���C�=�+?�t�������^���G��V}�gx��c������{=��3goML�!�+�6K	��7zu��W��u�J��E�~���S*��C9��E=7�M��W�|��;^��TQ �O���%���Ό��U�P��<��������������..�ȋ�C��=#��qwI��	�&����O_a��i��|��n|/�]��x�񼓵�>�$����#]߃�_�(���}���P%��[��5����k/�侗����;����,�F�D�+��^��_'ݸ��}��L�~���X;��gh�����z4������n]#Lcǽ��uΏ����[	�/]�/-b֍/cؿ����t���C�o�8*e����o���xT����k��Ow���gV���<����^��9
.���@��|9��/>8�&��v{q7�/������?^/�7ux�2�S���k�V�o*��b~՗=����O]}?J��u��E��(��~������?���ק��]��Kݲ�zk�׿�7��^���^y�xK����>����;��;.{0��WO�_��?�+�8x�Nv\�>����P��gT�9�Cٿ�sKWE��DJ��_���}����=i��~R�B�/돷ſ�wK���Zv;_�-��v��˫ ����(�Sc�u�����C����Hı}h�a����ު�Q��ܗ�b�`��]',�mv _^�X�(x�AYJc��*�-:P�J#�����׹ǣ�ґfe����)q��A�'��c����5$7X%�aw[�q$�P#�[��h;3������Ԅj�Q~�탬�=ݲD���^�	�3#��WuO���|F�3�35�ȣ�;s��c�hC������m!5�5�Y�7'��b}�KΗ�LN_u�t�l�*h��o�O�Fq�	i�ʳ��ԅ�M�F�ۏ�� ��-�\<�:,5]h>ȉ�Nł��z�0���0�mI�����8'&r�B���KP7�X"^5���:�aR�!�P���b�B�j�xD�:��&�dR����u�W�	4��<�� |-����b��=Rq����r*`���-(�^��8�8#�#6��0��cU\wjN�i�e�`\T���bXf-�@PO��: �N_���ǵDL~�۸�5���tg��M�R����B9	)�]X��N��2jp;���Y��f\����&����A��J 9�8���j(��C.�\�p��<�qLB#X<l��w*���9�o�C)��5�,��g	�<�DvH��!����D�9p�v���]:���дC�:�FF��"��4Kj��p�_Kk��ӝ�ok	��A�l�VFL�;`�������N��..�;����L/涸Yjp�sѴ�Y1�*�9��-D�h����0�*~~3P l/!r�S�Ǚ���p�(d�P��x��dN��v6�b���4Γ��7c��1�;��<O4��V�m�t�d��F�/���x1~{n2)�9kD��kôRD�3(C���Ñ���3��K�Cq��M��j�)�@�	C∳"��ћ!B�@��kBǩ�]
@tb�rS�F�,"	D���l�%%�8� �`�3����9U0>�w�i:n��.��ƸAo㱍N��7��L�����ˣ$��l�
�*4���ay�o� �4�Iy`�-�����b,�g��<�ڵ�7
��_2(4�l&����>��Ǎ��\��� �G� �H]B����%��Z���M���5/؛�1Н9)s���^�G($U�@p2�U���� ICǌt�7,��aN�o	m��ʐ�i_�.Y�v@�{�<�U� �KK�ȼU���
tn��G9���)h�wC����q�E+ĸ[��RT�Q�0G�5 n�qV��V�;��ò�'M25�e�K5�/��҈6�@O0G
�w�<�*��o_7�k}4����N�*��Ru�Q�چ>`�f᥵�:Zu9"��l�&�(40�}�2��D� �,��N��#�!�q�V<3F�y��X���/bt l者5l ���ڴ�R�㠕0�i��7��t������zF�0�)�O�y8���L�OZ�oIX��j��u6����|�qhUl��3�����s򚑲��[���n�� |:��c�m��vY���J@(�(`]����Ivc��n��8j���֜0<IB���~j� �M&c�F� S�y���e�r�Y��0������{~2���w��Xg�!�;|J؂,0ʬ�t4y�g�UZ�/f�Fv3�TE��x��&ϖ%*��-Z�:�@#T�r����-�7�4bu#���7j����  
*(��f�;Ľ�1Yv��>Cq弥)�)>�Ag����q^c��4�s$��&�VM�`Nl]�tbJCIKO�\���ɔt��3k�U��	6������\[���tU��81F!Us��v2N�jy�\Z5����ֿ&L/�$윬�@����Y�I%ȟr�>��l�Kt�ٓ�Y�L����[zȝf�gy#�˜�N���;FCn�;�F�.L<b����������5�"HC�T4�JV�yX:UӼ|B����VYⵑ���0�ڍ�t"��=w@��U�;	���=�A��`\bn*���Ҥ\k��ǎ�yy�d��ҤM�c�/��?����4����-��!��-_I6�@V嶤�H���Yӕ�Jdi�0�s�P��͜D}���+Q0�������v�YVX������������*�|��&���\�~!M�G3#���<�0���;�٫4�OpO�ry��^�.Kg�ɤn�D�8��B
F�~×	?i�Sh�G$�$�@�n�9b!�*4��7d�t ���Wu#c'A�⼠Zv�k�!�g��%JX�59���d�$qd�\�t[`�f���f��X�%�!F`��t��J2 ��89@(�R�(@�^W��H'a�i�msP�c\�V�A�)%�������}8fE��P�6B���a�@���܌�Y������D��0C����@�e(%@1Y#���a]c�*h�M�ǈ�m-��|ǮQ��������1 �C�qc�;*���q冡jU�o.��sږ�1�n6�Y8.���;jq�L6	���y�ЅV��kϚ!ԩSZܙ �f�I��Yd��L���k����)
#'Q�������㫂-`[��u;i�DA��Q0�K;,�q@ݠ��������XRnƱq� ��Y���?�M�����.&0du,m�������ǄbFXTA�Tflg&��,��W@h�Z���9r`G9f�
ƒp���1��o������)��>T�R�]�lj�݃o�JBܹ��C*��Q���w�M��;�y�k��^W5P��4���t�2���_\+E*^Y���8p/V�y�a�6Kw�h��v��H9pc���R�c���'[L�@�9��-1������Mn����!�k���s��ݛ�r>��j;����(Kr=�vG�^ :��dG��l�Xm���!mx��#�d�.!k]3�v�y�������{h5D��FL.��������G-�=���d�����
)�ɀK�
o�Q>��ia�2`#��;���L�3�m�Uh����1�����%$G����N��m�Q���@���R��*c���\�����	Xn�r�e�8[�a��D����A��v�K)G�����r�m�R�+}@/�Y�Wk����KB7��� <���F�6Uc]Az�bQ(�&/���ON�j8f;��������1D$y}*���pa1X�\�elĠ��!� 9U��N���ëxnQL��:zH�D�H�ą����v�zZv��,[AVS��
��Շ��Gh:h��g�C���p�	����g}>�n�k-6e?X�]�I��a�S���`4q�0.�Q�51+�Q�� �`��R�a��;Pd����O��
�d������(����X9Z���Ϟ<6���e������+?�����7~ �/��~��t�@���,�1�����q���X�Đ=����¶+/�VV9�Hݥ��r׹�@C�]E�`�����'J(�9�LW!k��E-3��>O��2$��la�L�F͓-]!B�/u�ܢ�+v�b"U�Y�������r\���DǂC5ç]�G�Y��фI��;vcL�(�,q32���I��(\�����a��@�� @�՞I��iF�CE�7��:<��t�A<&̏�l'�ϲ��g>��TaS7\�O�W=".�$�S�Z"oZa�j�.!"*��N����<h���.��r���ߑ/���h����Ks��8E�9�ԩ�Ô	TjT����	��	;�x�H��㝶�g���lȳ�����A�u�Cg*���T���/�
�Z�\N;�b���U����(��'�>���4<| ���<���!zQwP��S�5!&x=a{�_��J��DQ���_Dn+���� ��Y+�P��:�QH�� kx�ۚG���c��B�̳��6���|��U�!-�o�T�D=� 5�O���zr�� d��$�|�Bs�z��)a���պ6;X<d��Mf D뉐l��qJ��WT�}���!ɴ�k�F��+�f�O4�d5Sf���i��Y�aƂkWkn��Ԅ���nF����֝���X����ό+K�1pvam�ܻR�1ZȔG��YAF΅�pX�p`����0si6w�`r�h%��Ȭ�4s[�mw��x�N�	Ԙ#pZ<12~���[^)k4ڢ�b���v��l$��:"X��B4;��ߺM��I�!�	"��H�yo<n&���fW3<u�وR3��,Fh'� �k9��s̫䓖��A�*o�� #�s��L�wL�g�=�et�zE;q@�`7y�}đÉi�t���'��a1�gӰSL��y��q��0���4�	9���J��0dQ�,0B��<�56��31�Rb��MpB`p��G����a�P:�<*��%��\)�H"};�4-��{H���_�F2}�����-�I ��w�eBI֫�E��!½�<?� �L��x\= �nx� ��l���}=kz���h[q]�	��K��b�F�Z�#q�0Y ���r��N=�vv_L]b\p�[6�8�8�!n���*�xTF.��d�#b���l����μ�%��2�W'd�mtA��1�]���$@��H�
B����m�_��H8o����I�b���|��HI\�__Ȳ9v�ue�/9gR(6��3�U\8��C�4�O  �&[ Q&ӭ >�(���be��g(�
a*��J������:�J���Vr\-�4[��k����3Կl�m��k�M��V5���Ul�pd���HFI��e9r߳�)�cl�ʊ���&4?�zV�49���׬/F�Iwm��r�a�rL52WA������*i�p�4��т���NI��̮g�M��r�=�2�������e)(Լ�9��Wl�>��K*��z�T �Ft�	p�^y�aH�6�WK��Ҧ��o8�%��F�p%GNQy5J
�T)�08�b�npY�	l(��Y���վ�n���&���Q��mCء� ��WO�S�f��5C��ΣaW��eȋmk<^2W_��82G�	����Vbشl��1��e��؋��*a��%�`��,sOpH�v��R�8��5Fǖ��$�\�"��ڷS�Me!!����$}�6٨5	���,��BDU��T�o��Ƣ!IՈ�B
`"5Ff+Qe��:�b���p(E�Z=	&kt(a��E��zW�q<�#�����+t�Y�^���ՆvƲԊK��#�I���VE��� �7���=AY����vl�O�K�kVd9P��m�tw輛}��i�:y$�m��k�"�D\�\35�<x^��6-^Y�A��V�o�*Ϋ�v�UH���Չ��{�T��p�,�o��di��R�k�чu�Z(MI�j�
��^,���4�*�/�g�!&ظ��Ȼ��մs���<���_��.��C�X�ؐz�8�V�t�G�Cs�FF=�����L��Ξ��<1�3ee����uf�%s�a_s�3�cLSF�&���yP�Fj�q��FS�J�|���=����t�Sq)b��#7����[ȁ�3i�"��������f�]@K=� ����3NWV lj�I,,+��:��7D�$�k&�$s��.-��	��@L�a-�d����@��F��-�Um8C~=bFf�6�Bs���W���ߠL�/B%�� Z��37���3�^̀����4�,h}� ���l�g�6PC� | ���e��`^�u�r��`��śW���M���&ѱ�q5�8�VЌbK�14k�{�)t&nE�ɪ���h��p$m����?��͖a f���va��d����FS�j��CEd&Ɗ_Im�:(YG�47��B�|Ej�v&Qr݋ڀt�1�r�a2N���c;�:zi�~�Ő�5w��"W+��C�����X���m=�o�Fqi衛Sz`��M��. ܗ�Pa]�D��I:8V=�'�4�s����FS�#�[�<'b!$M�E{9U����a�Z����"Q%�7W"���]��[(2��C9�6q�i��MWP�y!׊���+� �J�R�]��&p�5p��o��f�#:�Z��Y��0��h���l�ow�3%J�:�ʉ0<=�h�M^��bϠ��Nv(ͺ�[\�C��m§�K�ήm�u��'C�����ݍF��LCϐZ���y�������Ky�x �ΦBΘ����~�|tnħl+	� Cm.�e�߲��m��
���'�2���^vr+J�A�7������;�<�	� l��_��D��~��묚u>����7`�����iK;���	�����9ǆ@"��յ�XAݰ��6�Zte�(�v]\k��"�C��@���x�?����DT1P��nbM���&��]D� ��%��,��!)��f�1c�������� ����H�m,H_Ւ��ܙ�u$+,"-&\-K6�$���#S�?C[�H/�B%CQ�sh��.J�0�˕ٰ��+@��fa���(��0��d�-b��0.���Y�����K�u�~&�*��S�BA��S������а�-���el�H4�h��&~�1O*V�)*
�_.>Urd�.�T~yv.��v.V��]s��b��2Ꙣ�jG��u�c����6÷�3Ͳnƣ�|SQ|�y �! c'���y�=q
8҂��%uզ�B'�$�'�.��"x-�X��9�N���.\��?
9�MA?U"`9�
1��'��������JE���d���~%�W�H��=p��3+�Jy�Y.w��e��s�������*|>^���z帞���6ӕ�[��O���$t�U�U|�W|�u�-1/o�/�鈷`����:��6`�/�b�>����<�;���SV�O�&~�۳� ��BzY�����I�e}#nK��D���+ޒ}}=���"�z#!]՗�`�Otg� ��P ��߷W��a�]�oȬ/��T�?=��נ���R�ik���Y�	Z']}c�W:��W����ꆻ{H���(m��A���_�+}�M���j�����g?�ع�]������&������o�z|�f{�O/	�.T����;���@O-vu�׊�SDY[��̈́_M��.>�����dر�枧��{�\�Ԟ~
=W�vs��$��43����K����߳݁M𕺾k��7��� W�#��;��]���,#@�`�����������:�[p�7��w��"�O�|m��q�zmw �y:ɽ���\0=�2��kz@>3�R»z(��k/1��6﶑���������6�(f't����{����ܝd�Gꋬ�R�1�zt�� �ܵ�ҦA�g=*�;����)(�诒_lť>�'��c���O9��\��n�0�㏨�/c���҆�~�҇��o���1:�3�>����N��ϟB>S�=�k!��>;�Ë�s��>����釧�YY��|��d�{����m���'��G(�)�D�毮(�[�x��4�_��C�
�C?�/���s����X�R�_�2�H.Su�#+��r{��	�f/������I�}�����������<�uq'm��h��Z8e��eW����z�Y8��S�G�_o���~
?6�j�����������V�W��_>�4/��+o`"�٫{m���F����V� ob�74�{۝�ީ�ua�s>�ow�{/_��m?�ߤ�o������"� 
{����Z�k�_���M�7�rɮ�k�#�����H?Fg��t��j�6L�T�cW-���,�ĺ�4����/Y(�ݽ8-�7�t�W�����~62_�M~�灍t���u������Ww�s�	�G9~|�=>��Pny߷�g���ꝻSxOB���R]�f������NW����Tl����T��^g�ګ����ry/�A56�zs����0|WR�o������]vC�^-�����*3�3��c�;p?�|�'g�C:�����:7�'��+}���ǟrq�!��_��~�~y��rb=�����o�E�J�}���M�
��?������z흊�Q��=�꛷���j�J'�Q��z5�D�y�������O�^�R�N����Q��}9�1jJ�l]e-;��
�y����3�&��mc�z�z����ˢ�o`�������J}*u]����	�{}���$�����4����	�G|^��w�lˏ,��h=*�)�����&���b������m� �lg�y��`����R����7�(����Oe �7��~�oZ����@��v3R(����C|�<xz�Á<�~e���աc_z�}�ޏ]�q`���ܿ���c֓�z���r���ѽG;'���O?ό����%V~mKR�tH�O�<�9K�ؓ���	�W�w��޺�&g) ���)?R�<� x0�������rK5'���;I�b�յ�_�{����i70�w?M�7I�=̞�]Im1#g��[��2oѶ}�i���dm4�_Im8�n��� �+s��������^�_��|^�{����u���F�D~?}��r�kxD�G�����sx���f���͐慧�yw���m��7��q����ܑ(���N>�/O�^d#�7%�ܙ�omF��� ����1}����M��LP��^+/'���*��##��%*�/�`�7;�ϋ�z�v:�_�,����i�i(�HU2���`^��^�n��}��%���7��w�4�O�����>ɚ��������5�C9�7��d�5��W��d�\��4�W_K��������׽:\�����Pr��45�F"����beP�_"3�M���;{m�:�g��y0oU������:�|��g�R5.���H�u���Jv,����]��m���O��-�/��a�Ы����z_d������{	�{;�|���۰�o?��[�3{�Q^X-3�0������#��ALJ���>��9Ǯ�����j�bĲ�Pj�pc �0d��W&�d>H���kc���j������m��]��:�s��"�d��9��k`�hV�G��+p䁰F���D����6�~���e3�K�5���3YI�c�[2[�37�,vK��sX����*�3:��;���ݠ��[%�C�
�����`���թ]%�<#�U��&�kE")�<��!󐥸"6�g���C�`xÎ�8�d�J�ˀ�g�0����	�Ϭ$�����̪���o��3a��Mҥy�`����(|i��6	��y%�6�=ndKkv  �1Q5|H�� h������P!�{&Ńm�r
KZbo+'���
�B@r��5�r|�0M�se��A\��b�B{�Y�T��D[k�\2�4��FSI!�A������p�}�	�2Q<�ȩ[v��8�&�-�K�a�&\�*p�!��7v�#����-{�kA�R����N���cl6o0[�8��xL<�E��TX�Q�����e��Y0�2��5�C"ˇf���؍yrD�
�b�_d�Cɟa�/�ڗ�RU��D���pibt���G�yP�*�Â#H����p��L!��h�m
#[~+�َC���a3vQ���PON/�Y0���R~�l�"w3O�*�'da��L!��l^��(K��'���`��n��3�z�,tJC�f;f\h��:���U�ig����ቔ����m���#_h�d/T'��`�DWFC%�C��/:>I�ҞQa5��R���fkW״(|�m����qP^�H�SK �+�MU��f�#'O�M�����ܱ�k�2���V��ȕ(7Gj]s�
���g�v Ctj̕��&gr�V`��Q"�2[(�*���y���`1Ȕ����!~�yb�T��0���]M^X�]�9��"�}-[	��"��Ȱ�S�OY�%L�����(g{E����Y,,b�6A�x9>+��Ob7T�4�W���jc����Đc�_k�:��af�8����1�;����8ڍv,WiS+G0�$�$0�ˬsc���IY&]�� '��M]s��2�J.�6v��:�VB���`�D��j���w����TឩlE"��3)�gT�e\�x�{�--�k� Ɣ��v{�ӱ��C�ׂ��gI���R�HKq��nc#
[���S�F�9NE�py>����C�%��<^%���or���0�tvE��4/s'��� <�aN�8F3��܌-˲��bM,�f�U-%!��t��(��X���7�_4��kq���e�o�)TLb�~� )�0��5O�h�7�,�@a�\�0%�gX�� [G�fF�a�}��@�����t����J�%�Jc�e}wΤc�Z�ɵ!mM��m��%'�|�FR,޹��qc ֒�䷴풼���	Ѵa�10��!����mNR{�4�Ya��A��#xf��UT�}���D�uw_�����T���z�PV`�xQo����GѶ�/2��.��>�3��e]LȊ��x�F�ċ#�5�Ot�u�Y�a����� W�^�v/��A��,�&��n