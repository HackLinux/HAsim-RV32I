+�Z5>Y#�r�������3�2�f6�O�gPQvVh��a���<[��R~�H�ht�$Ɯ�?	_�Myi������c��'����ۅ}h�'h��5J�s�{������ǁiᆕ�4���F����G�Q�{��}���E�j�_S��ՁM��c�#(�#�u�Pʌ��e�+5��w%M���5 ~؟NJ=&���+��MY�IG�ڙ�Ɲ������폣��_z�)Oґ�Vj�J*n��Q+�91�*�(� i�Ww,��@X������~������ֶ |])�.����؝��h5%	}���z��Q����/��w?=&��\��k6H�A���X����W�,���A���DuS���67��A������kD=��5p��`�`���<�vw�ͷn�
�W�iշ���d�J�����iFs	q��y�>�'�Kf�j�Dx�7��1X�yp�E��3����:�~2�W��~�q�_-yY��ٶ��}f��d�߮M<���~��N�ߦ}���uy��][���/��.;�m.ZƏ��H�}��y���Tg?�"�����XDZs�c���cݖ�>	�+��Ɵ�����l_�S�5���>���Q||K��у�R�����сã��O������W����Ӗ67�W���@T  E�D-�{��Z=���"g�0=�q1c��a7h9
�l)�(@J�
�t�Yc�n5��/e�o�2� ը�;�������Z� (�!�V�;{j�!N�6�P�\Iw�)hb����Ɯ{�td���W�����{{+h��1"���^U�Yls�t�͓�K5���`��ΠBk����ʝ7yN�X0	R��'�ܣ���E�iRP-T�%�+%�eX��^�t����_[�Γ>x�uL񷿡������En���.=�~�5cPt�"�V�<�v�
�B��ygzczk�F����!�e�Je�kM]n�3Y���\̎�u�_��jx��0����/ŗuH�^�)'{n�ȁ�M�4&a3�M�#hf�{�~r��?�e��A�R32?���`|���w/���ԏq���e����Uwӽ��e2���WO��ͺ�D���"���{kE��7�-�����	��}�+G�=�{@�81���_M��dM-}��?���g����[P"�MaI�
`��(3���B,�;�J|G!�?��T�-��;
�[8���`���ȟI�^��Q
<�O}�����=��qz{� @h�1u�]�����ny�����=����[xT}{�_��B��|��������9g��<�L���������ʯh4環��f��1e��U��BCvM�l['r"�W�=b�l�ϸՓ��P�hV�b��G��Uϰχ8�j������1w;���L���_���Ch�Ѥ��1�[^�����������e�r�n�yjDG��@���|���"������9���y_�|�;#*^Q����!!����h\O�_sƢX�
�a�h�m'#���^p�0�] ���.��xc";y���	�U��?\�N�>>:���:84���133�E�%j��D�H�`E�-8�`� u��`E�%:� ��qr`A�8�����s��Ć62p��
�/h D��k �)G*CY����,Xp`�
�6��%:� ��q|��D�-8``��o�J��ą�3 <��D�%X ā��j�t�̺�*�V@���Y��D�&ؙh6��0���#��t2�Ȁ���d���O@ 40�̾��4����2Pj�\�P�Lp��J :��:<ܾ�,<t� 1����