�y�q�_=���m��XCXׇS�s�;_+��<Rg�ZM�9�P�P$HA���qk������x�A��@�U���) e�	7�ۗ~�z��'�s��bp��zz<�J�*�p:)Ň��!�]�7
�}�;�\Z�Þ��b�yO���>�1�����*Y�J!�8�ҳڟ.g��9�O)�2�%I6���1�.��b��Gf 2z�����1�vU1�R ۵Hl���z�ϧ�w0cT�G�Yf��r�6w+W��b`���z�<hHi��8��v�y7o����>^�?{���;7j���_" �V�6/j�ze�j��p\ȳ��M���T�%O�W���1$�	` .]�~oôԮ��p~��s���ծVM��]9�Y������K+Q�.�z�TE��
V=����`p�
,�x�<�H	�J�@���@�������ԒX� X=4y�%=�c8c����M\�p��^�ٝ�r��RͿ'�ԑQi�Mġ8$�Di R'P�@f��ƈB� 'coc e^��n lRa}�p�^'{���ڭ�!�>OO�����bp�
ܻx�0�H	Pn��DH��~��]d� �x�	`�V0�(Ȕ��J���S��gM���o�����H�܁%6�:��V����n[ ����<��(��S���d��Y����4����ڝ���P�U��G��~}���PV���f�H���bB���b`�=x�$�\��
���pw񔮨۲�䑭��Tg	[r�
����T�<6��_wҊ8N6MнH��(Ȝ@�_�#���߬Р����f0������pp�`��GÇ�*��N/v�����j�����׷�Y^�F۔eHߌ�X�g6�J(��``�	��xzIH&��J )Q�"����͐���ws�i[t�e��4��J^��YwWm~(�0�����iE���VS���|���!�6�g�|.�o������~�L���	;�������Q��� ȹ9&ſ|X�]����Di|���bp�
��x�<lH	
�l8�q���嶯7���&Fn�TLLJi����)l,�cm[L���bm��#��r�˂R��&���Gz�'�{���B�>� �ǔ��]>��`T�j�r�0�Ӛ1𗸥
[��~F���u�O�8���#�_��bp�\�zlH	!�p(�q�X���$BK�̌8r��7"xfJE�0�5�rKw���)Z���H���G�z��Cm���B�c�ɸ����~���e�)�?2���m�(�;��������TS-#�N����47�RM��Q��߹H���U�C[oO��F��b`��}|�%(\��^�p�9��mj���������Wv���^gK'����Me���-4ONf�G��F`���� Ga����g�����;+/��O.����V�r���g��Ի	 �|Ej�&Ŷ `��yB����sz�E!A a*ʜ��``�Mszz �\������p ]����䯑"����kĻ/~�4 +U)(��]���ƃ! ���#9��<�+%�D	":�,A1�VHkO��X���^En����s�k�8�	N�H�\�@%9��}X��q��FI��:=�ȩ�XYU����bpo�z#HȆ� FH����9� +z?9���*9ݺ5Ԝw3�Te����aSEM.��F)��FM؈1�S�}Cz�o�4�S��oS)����j�D>eT;��� �R�B7�e�J6��)���یi	̪T�')�w���BCqID��bp�	�z�$�H�*�p��I#�	*�2�^�NKI.����EJ�$gXˎM��~_k��n�0�s3�_v�����%�b֤���5�4�s'QT�cv6�eX�A3��,Fl�U�F܌=4켆J�c�kC�e�����_�������bp��z�%	H	�Z� F({8�&+L=`-��0�;���S	�@���9L����Fڈ��};���������n�J�$����Ӵ ��'�f��z��Q����1]BCq��0��R6��!Gr�u9n�
k�b���^�|�V���s�k�|���`p��cz�1e\	1�pJq$�EA���B��AI�%5@�y����z*>=�j��I�ϣG��Ҁ,0RV�o�q�p���!����Ｎ�fEY�W^��Z�����ԋ��N���ߎU֬�qPU��F۸�e�!��a�31s��D �̍��b`�
��z%	HAV���D�������Ej\U�(�%����j����}���{��S�&��&���!����h,�E�&�@����ȧ3��J��b������4�a+�����䖿�q��(#LR�kՁb(�).#kYi�FfJ�c0�)9����bp�
��z� �H	�� Jq�� �̓���m>)mlR��*�eF���I��e-I�T/|�Qۿ�I	u�v��_�Z�F�I����C�+��:�_%�;3?[�򫔈$�"�f��J4�Z�nH�j��h�p�9��������E�m���|����BZP����bp�h�x{%	H
)� 0�q�5�z�l��$)�ŅD�CB���u�/�]��=�I����{|?�U"�(��	$*}{� �E;��������'z��1���Y������V��ې���b�/��d����0�#q��](�}���JM��A�2D���`p��a|�%e\���Dq���8B݋D��Q(��!r��ZM�<����u5v�����}���{sU�(�椲�5�SB,M6.�
0 ��O��fu1_Ԍ���o3�=fiQ������]���Ϳ�_��~<�} eZ�Hܰ	��&�>[�T�|��b`�-gz�1'\²�����c��Pt�#��jQ��K�o�$��)<ʍ<H����TBD�4%c�hwS�e��WnQʷ*=@�����a�"�;�T#321�����_\��uyW�ވ����[���r&ɿ��]��o�gz��Z��ܰ(ƇlR�����b`�	��|�,�Hڲ����zW���YRw��Xy�Q���{�E��厮<:\bb($+�-E� �o���[?����eդ�c J����G5.V嵟Z�$�@7����o�h������]��Ĉ*�^���
B0Dz+SG�3��GH���B�?��`p�4�x�<�H��pIDqP��ޫS��
m����#�I$����Ĥ�Z�P����]�wwV)����D�"LA؛`�!]ߊ��~
�E2$Z{�J#4'AV��P�Z��`d#7����w�*M��_���Sa����'��q�r*����bp�
�|�$iH؆� �H3K�Ш8 �ҧH�i#�L$r���z�jV�m�O�ҿ����F��kh{��[-[�+0��a�`2��)���Y�9�W9:���D�;�,�^
��V��Nݴ��Ң��%eM%?�-W%{�l>G+!2k��Vu*rr��bp�Esx{1'\	AN�X	Ɛ��
eA�
p
`�X,h�#ˊB� q!����q�Q�Wwc�*ݨȮ�Ov�gjgM���ѫ����ʹ�)i`�۠@U��e�F���8�����X��<���y�am�KԄ���' U�<�_�����f��Z�����֛�u����b`�9qvz1'\1F��0����Cg�m�`E)�i���[�H�������Lۚ(��]�D@*�4�����ݠ����}{{u�i����P�ʣ����L��;���l�I��Oذ �U��$,����m�Wr�H��T,�Y�B73�{��8v��`p�	�z�<iH`2�T�?���@�0ryP����HO;!�����{����?i'7�c�ևOX*jN�irn�s���lQŪ�}Rn�+�EDq�~?���$�܃U�A�b�>p��Z��$��v+������n�ƒRT��t�����
����ALk��bp��zz fZ���\DL�H�C�j0n
�z�) ��J�?bI�>k�yF��	L� r���(��u��f�qw��K/����ؑ܏'i��Z>_�*�F����A�-�93h�b�.�a��M�n�@e�Q�ܯ��J�3}c��թ��V(���b`��w~�=\�Hf��FHU��q���KS�}
�����h���#�nb��O����Nk,=��w�ti��r�͐���6լmHXeF�'C�D]���  bI�%��*t��W(��NrT�c�n�׎F��	V��8Ľ�g��ŗV�A D����bp�	��|�<(H	R�D(aI��Y�a�����GuT���_#3�M��a|�U�E"�J��
*C�;Ub�P��O&��8�ݴL�ň(*%$(@(��@���v���6ɇx�� �F��n �.$�����\����fh,8S�g�T��`p��v�<iH�
� 0  ��i��)�J�s��!=Mp��
U���UN�r�+5պ�s��M��w=`�g�q- 3ֵ���L�/�I�����%x�$<�M�Lbm��L�Xv�_(��n7$�����Ҹ�?��:��!�NTGq��(������T��bp�8�t�<iH��r�l(DH(br���� ����� �k��?�]b�t���麄���2.�j}�����iU8�����4I,K"m�g�f����%�{d�n�;���9�u�jw���j���+��W�ZZ�l����Ƨ2����y��bp�c|,h\	�"� D�����M�<e�ۢb0�J8I�h1ţG"?c9�fER�V5��K���݌�z�-�D3�1��S����da��`�B�"*U�c��D�گ�@���=EX<��W����z��:�fJDj��ݟsMy7L���?uj��bp�=Wxz<�\�x&�p0F �,�Y�u��tMHFQP��Le+Tȓ�)��k�����[�m�/Uo��˴���M�U�(��Ȯ���]��H���@�uU��b��p���Ɗ�Hh�h�u�v�"wC�4�M�5Q�Y�le���ZB�����`p�ecrj<�\��T�H�3l�"���5��\
�<8.�0��\���(1�8�ɳ�F�I&-Z��n�[��a!��-��K6/��Z�[@4!G �V���<�7J�c��S.j���g�{v���q���Lץ�4�@`v�-
�� Kӹq�5���bp�P�pj=)H���0Fqe(�,cf�3�����������n^;�J�/��ӫ��2�lX<n�M� 29%,i0�i���ΟXqh\��/����o��/ЕE��n��C{�Ǵ�6%����63�[5�'9qx���H NP-0B��i�uS��bp��Ktz<�Z� 
�  ��"�v##1Ȉ�ʗ*��+�����t���E�8�Ue�qJRe