�m��W�wqF5���;7�S�-�
r��yR`��;��M&�E��e���d��9�����È\N�.>/H��I�c�.Qti,�.6�y�;�����=�1�v�-��@ǫȮ��V���c��e�T���la<tڭ����>�5� �\i���CG��8>)���q���h�7`E��sĝz%�K�o'=ʱ��e*m\g�A�Bt�В鶿����oF��.���.��ݩe��m�O�������Zd~�\�!=+�zn1I���j�.�
v%Q-p�,�-�ɺ�/J�-g#z�k�҈�׳G��2X��i(�*L�����d�&���4d�I�5ɦ&]����ХǭkHLj���f��Z��+3��(�묢ýة�U*��������U-D#G�BxMg�!3B��!V�JA_��o�|��5ܛZ�"�Ub���)�0��5�Ck������e�4W�������Xw�D�}��v�h9Z&D�g�#uh�6��\�[?ـ���!�Q�4��|o	����0f���1�b�
[�}��N�U�a�l�d��9�~�k�7��ߜV�]N+��"�U�o8�~õn�+��쯜Vp�rZ����i��+�<ѯ�g��^%��p������o����~ÿ��B���o���~ŞI��i���WN+T��p����i���<� ����o��pdQ��ӊ�7�Ǳ�+��7����7�o��W��rZq���߼QZ�A[���B��?ȿ� @�������	�_��ef���������<�����^zq�k{�X�A��l�R���r/�c$ᢈe��<�$o�g�%U��:���5�j�j�kR�����!�=�P�+w���½��sތ\w#,���1�}�ב������Z[���|����%���K��\����w�t�����{�3���6��w���|K���[�PC�����֤��ǃ��c��D��q��lU0�v+��@�T��J@�VB�Đ�5?Bp"�,Q�T��w?w[&�=�@V-X�Bi=�>\���g���֤L����W��l�������5��;ti"X<���?h�:�Jw�/-��9HB�z����<T�S�.�9,�[�N\ogH)�iJ�/�I��� g�rC��I]��N
>s�Q��CmnV�8&�
.�Y�`0o����`��g"	X��qE��m�K����'�z���r+A@[Rb�)C*��x�h�}�vG��X"��2ʄ�J�Z�k�Y>|�$˖����n�(,�L\�o�r:���SV:%�F�3�������}���2:{��V�La��ex�q��t�r�|m�*��x*4( &G��r���҉����3�7�}N]�,z�j���;�߈F�W�gy�
R�}��}+�E�[Z,�,`UA]�9�"mҁ�X�J!���X�ڴ��� ���.u$-FY�`�ʀ����tv�J��>�H��1�@�a�d|ٮ��H&�^$�[��/�$��4�o1��e���&J�ֲU���-9��
w�0�B�+�A��K�@:'�᥯/�
��w7�W�"��� �E�TS���_�ف��� ��q�d�_B�U0��7��t���sp�56��òvIx�X��{Nd@M#2ow {�(1��Zr��y�;g�8g�v p�,:jz�F�%���$
����L!�8D����#H?��t��������Qf�=�q~#��΀��6eΐ1�)m���ufix]���g���Ż"�z��oc@�0)HJ���:I��>���'c�k5L
���,��=��!,������S�����^�7�	~�8��������u�����ί�] �9�B޹!9^�������Ax���jP�Q�Ӗ�Ry���s��1K(C�쌯"��UF�Eӛ�H��hPsp����[�RĻ\�%��|xqS	����R
c�C�#�'�7�NA��bǝ,!����[�w|�T���np��3zd��dX��kV��
���?�9l�y��{�=��7�HG-B�ie�fV-��Zt���7�+C+����#�ݺ�
4�tYi@X�3��"�;�����j��}/�P�O��N�mzR[#j�n�=�k[��'�,`-�[ɔ8�,;���i�|���Xjd7�-�
(朇,^P�`�6ݽ�ĝ�;�{�	onz�� �m>!�8Q��d�w��BLQ͸�s7��>��.=@��M�$yV՛�[T�{g���fW�J%/Z�	�Q<�X����b(��g"�!Դ��W���b���C�p����F{�.�a�
�o��ŋԋG4.+�ËaF�F�5:��X)fX�]t��)Ԩ��Ʒ��O�a>�l\s�)�XUF�A���NJ�������sܣ�6�*�56D��UyiE����n ys��B�������g#�A��ot��Y�=#�G��O���&��O�׾��D�#+b�mO�&' {K��&�嶍�H��NA��0�͋�2�яqX  (9@i����x
�> T��Γ��O�e��ހP>}��d�<�Oz�>�?��̋'3����dN�/=��O�'>������)|���'V�3Ƹ����{�\�j��-�r��{�15�^��{��x����7�o���{�/�s���y��5�s��E�s��kMs<Ut�&��.�*��bN3N��l~Ӷl�����{�% �su�,g�}��<M�mb$h�ɼ���h$o����
AV�j�0B}�9��x�`�`ص7q5��4���{�î��k��u�H�)�0��m�k:����g�h?���3\B\�S��(�ܬ9��{AU��^�S�cd����/Ǝn�㡔�܃����S���������+��%�V_�(�,���`��a��^���3����|�|���e�a�"Qt�^��z7�"e̥5[�?�~Z��6�A�x�%��&c��Rԃ��@�Sa��d +HB3i��q�}5�J^�Ko��V2���7�!���?�~?��u�o!��J|��h��,i�e-T�)�'���ǁ���n�	����E�|���I�$�wRm��������!ín!F)G�#vA��0��7��cE5��O�/�?�>�I����u:ZlCm��H?���!-K�~��f(uRP]���ўf��\[;ݴ��u�#ān�T�dm�۞Z/D��9k@s�9)�J��/n�%�;���|zM��=e��,���!á�WG��295�V�Sn��.�CmCɆ/2���[-?��^P4ݠIs3�U�׫2��_��Aю|�:�U9k>��<�H�M�6���Ğ�#��[@�}K R#��"���������Ǟ��]H)��V��Κ]�f��n�a�#��U,��77u�k�ɠ��I*�ë�%8�H\y��=����赜l�ENS�k��&��%V뙹Vi�Zb5+�d�`?\�y�D�>�ŷ����mM!~oB>�r�zZ���9t����NT0�^U��¨\�9]�_g����ݦ�7�`�_�}�yZ-t�*<k)rs�j���cd����b�h���a�A��lX#�}04Y&�e��an?Ƒ����e,*��/ru6w�#�i�ok���	F�S��_)�IZ7��hV���Q9�Q���qM��{�|��75%n��#���1�+>R�]}	�Qg���%�Č�BR!�:_e
B��$���bX���>Q}4H���y�aj���Ȑ�w✐X�s,ۓ��mkl���FJ,d%'�H��� ,���᯺�K �CK��tI�(j133333Z̲������Y�-��b����Y�sO{gwo������v�;-����(��2�dF���l'�tar�� +f(�i3�{�r;�8��Х@�@���Yl8����2P��� �����5U��n���ע(@{���9pF,��B~�_BF������Fq��ʥ	Ѥ(@��	�P)�2�v�g=��^���!��Q��r�l
H���m�l����)��g&ɩ�'�J�f���vg�~A��7/	�[��wq�O{W\�t�v�.��D˙���Bqߵ���9X����t�M?aA� �݀�^!�Z�@�B���H��2��OYQ$I%�#����s������Cwbީ�0�XN~��c��i��qG��C���g�sj}92=k�p��|�_&5��m �n�u��I�XU�th���n�uz>.id�ˬ%��HvP�5�iT0�jhh������+�/n�<w�2*��z1�]�����!%R+~G>���:A��y�;��~\l}E�c�1~�𵣛k�A���s�B�'|�J�"Ymwm'+�ۋ�|mVS����áS�AJ�C�X��?q���1� �A����Xo����Ѹ\����-��:&�ڳ����@q��q.
��� ����k���1D�Ȩۛ�����dN��p#l9�\����.0:#�G���0�%�Yq��`<�uMăM��6{�{�L
���Tl��(��W�d�̑��.}���Mϡ���E��2>�ljO�4F6�����y����`��#�ÑS����s'�o�g�g؆t�U�JE�L��R��I*���&�F�IRDC��K<T��(��R�fV���Q� ��3�:�g���q�M�ܻkm�90��o��(���v]�wʡm�I	�<�*��ς����|�BJ�dRj����7~�-&mZ���7�FeY-�q��I�#�K�1#&?ЛG�����k����s����F־��E�e9��Y��C��5C�:2�J�=�٣7.�s�%�t���y�����JpڣW¦d�;��&�\o��)��A�tl����Ӎh��%褴y��O������Uv�_�u�S�Ǯ��.��8O�ݏ�>��Hoʯb8ݎmq��vn��}
<mdhp5M��7b�1o��.;k�'2�}l�B��{A�r�Qc��t$��!烟G|�^�Mk�|�0>KH��>@?F�l�٣s�����=h~��� �Y�K��Y������4O�^���������	Q�g�� �Dʿ�N�Ϯ�p���hm�"��cz�چ�6O���V�	U,nN'
�"=+$,=��"L���AFV�Ex	��@W�C� �k@�����0��T�	q��d��uv�����󩡵��}��t��tPy>y�"F�^"�a>e����L�ޱ>�d��즍W;�7��p�Zjc*����q��=ש���a���ic=�2!����n��ZaX��мvŘO-�m��:xR����d���Y�.��:B��`fA�[����_�����f�T����T���x��a�F��,�2���Cx�x��&'��*A_$��t�a!���t>�fF��/,����
�����P��i�`nY��i�M2�v:���(����o�/I�>���LS[�G|F�-V.�$��G�g����O�x	�N'F��H�\!��G�`�ƒr�½���9���٩D���A|*�x���߫��Cqf ����n��4>� ~-z ��qnR��o�w�� �8r�G�%�r���T�c"��tڌߧ�s��k�A�#LԾ,��{i��Gp	�%N��>��R1�����j�Y��]�%a��Ij-��߉���P@��m��^9�K��SO�-�FnUx�"�(��]�rd>(�G���|�CT�_�٩W��i�Ѳ�=�IJ`���P���9;�e��ONw:^e�A�=�v��3H�cp��hЧF,itpU/a�	�w,+�f'Y��bDp'P�U0�"N���B���]�w5�Szr��C�k4x��ń�0�7:��z�J|�t��a�����Y����ڥԚ���z7���m� �P��w�y9��Cs�����Ŗ��RX��qiY�lqRA&wך�w��9Cg�?{�f1gN��q�:���7�^�޼��:�vl��%�F0�n	���Z�Gn��E0��s�5|}d�LMG��`�V��if�&{�D]T�6]"�	&RS��f��z֜j���5��aev�RBT�ӞPOHK�������A��LM�ig=���"��99�E@��L�c5/ѩ,,�������'�[�ھ
b4 6�b^PM����Vƹ�~S�؅��"u<s�P(��!�v	�M�j1�l��,L:܁�z�QG�*%N��82�O����pB��t�/Nγ�'�!':z��W�Kg剖�g!9Sd:"����9v
;�Ļ��6��:(�jT�/]�E����H�}�g��lou5�[���� 5���	=>�I�be;�i�XB��t��z����7�d8j�)h�ʀA<�]2N�a?#�}�Gd�{�儚��6��-����+���mt�eA�=�٭�����_xU��E���2X�+S~�A�jo'�X��Jz$�Z(�M@]I$)ǵ�(���q��j�.*		�3Y}��x�n�@T��g����e���"�F����쵃
m��P�d���\�'f�k��{�ܪ�Q��U�x�Y�����{��X�\XY�o�����]=H�rm�X�^�Y����<�S/мw�
Զ��I��PNy�|�#��	�@ٳv;��FO���LO	z���e?h+I]�Rm�è�ew'����9,�J7�Pu鈆Ӷ蓊�6�?�4��iP����}͟��'��������U��,Iﰅ���^[򆇶�X�Cf#�3^͎�Q�'�K�����_c��js�@��F��/��
b��w�nY�J��H���m#�n�ǟ��:T���ﺱ��a��`i>��҄�ʼ�� �^�Ѱ�[8ɺ��g�;�l�}wq�xt �`�����uTF_t�+Z���H��K|��]d
��!rC߷ �o ��j�?B�ff��c�}6G����|�#.wi/�E����A~$�*/�� �e��t�\�7&W��+]��k�+�f��CVQ�����-����*��jG����/ٗ�g/�M�g:����<�OaZ���JB��Z(�a��LU�U���?d+0�$��\��}��ϯv¼
�����F�k���R�W��rÜ����}bi�=�x����7�8��揞����G�m�y�"x�[�F̷�q8&�|
���Y���$���x��,m�{��*���)y�P�#���*߻=��ݢ�Q4�D�Բn+]s��VPy�S���<*W�ʅ Q���P��j�����2� m���7�>���v�C�6@�]�bu��mzʚw�����k4G|Ұ�خgn��@ۘ"!ӂҠx՗�t��==���1������w�����úÿ�_��p��� r{�ἓ����������d�d�_����_ȃw����N�x�w���;mﴽ�3杶wL�;6~����a�����G������@~Ǿ�ؽ��ι���y����!�y���C���"}g�H߱9��t8�s`��(�o���lp�5�:����[�w�_�{��O��?�9�ٜ�����V毵2�,6����cdj�#S+�gm��ޢ�8�DT>S�v⿵9��{S��¡�>������A��>%[x�[�ƿ���Kk�o�1�6�<֛[ǉ�V4�zcbeYF3�59��Ol�͟���{mگ9q[g�3Q�k�T�k3���(�������9�?ɋ� !����������o��8��S��9�u~�:xp��N�>uκ��q�(F $]%����?�:��{���\�����7����o��U��pDQr�d��[2��R `� I>{�7Kl~B��(�k�<��ê%wg�8�f*�J��\1ŏh�H*��C�|����C/>�'�)?��{�{:�8�Zi�룞�k�k�Z�҃�_�2@3 ^v\��L� �z]#�y�z/��]X�zv�w��-���C�Bg��B>�ۥ�ᔑ��-��d��������	�����B�&U�DG��ԽmC��t	A��(�.	��y�}m��؎El��%���7��1Xm�u��$?Q6�o��$A1p�����(��9)�|0%2"�����A=�GL<#��	L��1���xX�.i����֣��˝"D-�T-KL����PQ�aYs�T��Ķ�@����%��8������Q�@���oa�O
�2=nx����8��m�R]�sP)�
]*lks]�K��Ӈ��PX��:��vǒ���t�6�s\' ��ŏ���'8�q����m�H�u��N`#ԭ�V����\p4���Ԙ"��)J����\E� D-G�yH��r��Z�wv��IY����2U,>{�+9� �j�6BJ�&~;w�C�Y1>�<O*mQ�HKS�#@Յ"?�nP��(7
d��o˙�����I]y<q�#��`�؛a�r��'��� ���������"Qy��"h_�'þ#OP��N�YoL�IB�&�'�I��CCmn� [���.���.K������/~VU��X0��c���FV������X��)X9�0I9K=2bs�.��
W)�r/�m'�ͧ��ӿѼ5�,n:DF�l�?[a���A�+^�_]|U6N�H_��)=@y,�崵�Y���!�e�8�}�4~�+%,r�Ҩ�?�J�*���!�Cu`[&���b@]�V,�6��C��4J��α����z�m��&Y����o�&���~���F�M����'Ă��YǱ7{wT+˥l��4
����[=cX��D:BR�9~OF]]uN�Uq<�uo�����T���Q���,�Wc������4�^���e5�\U&�.�]+w�OP�w�/ԩ��~���y�t�߱5�i��7����+ڌ��C|�5	��\8�ʸ����I��10�U�V��0�P���e��Ĩ��7wG�X��c�E뾪[�6#��Q��U_�t��_(�ʹ����%�j
��>�8������g�^��/�Ý�YZ�Y,=�K�t%	�� h�{�!¶�	�K���B3�Ep�!�k��*'U���I�8$4
�I��$5$�E"�0���P+N��M��uP;K�q���0/w��o�� ���C��X0 @ݯX��ϲ�k�C����/�����/4��T��{�~y�_5ï���~��5py����{ٯ˧_�گ���_�¯����i�߃�k����3*-a`���(0�yC���;T��bqe.=�Ѵ$����+f�W�⯘�?��a�����{����>� � ���x[!�c��@�r���!H�q�6$ 1�}��P���S  �XR�Y���ݏ-R���.���I)=-d�;��W���,���ed!��Jx������b��瞈4�s�������֢E�8\��k�������kOd���e�������d��E�|������^���oxlj��W�K{C0�P��Z5?X^d�F�*^��E`Ͽ�gc^Q�N]�qD�χ�V�~���%��,l�칒�$}�S��j��n��t��h3��9W+'��T<!��a�}5�G�y~C��# �
) �E�T:�hň���K�FBd���/D뭭0�m#�S��m��T��X�����<��Ks�f�/��ϴ�b�;I�--�B����O�e�������A#od��WL�_�����������5!������烸��ޠЇFB���9�������D�!9��NǛY� � ��SSy1킧���r-����Hs:3�#�&��|��G��۰7�)6��`k�ڗ����V[��]!�IÒ�KN>�<&�J��r�G_ـ��=9>������Z|�M��j	��\��_pcO�A2YFa��D񗹜���8���4�]���V�e�sd6]X������	u����K��XG���Z�t2��p�
�A]b�W�{)��5Z6�~1��<W���a�������6]P�F+�_�Z�yA��}7{@��gi�8�;��ߠJ��ƈ�'P���W�|S�j�� �y��x72>�(��f\܂�jjǞ��Oiz�,)WT`�ƫR�c%�-��O1/�)FW��Y����e��ͺq��N�v5+��:4���M0���t�u��!����"2�p���y�D�"��V��#H��J�Byh�'�B�2��#,�[;c�h$�����[\W����hb�Y>��J2ړ*6wTg�b�α���_}�����м?c�I�j�9�o����������� �t������[�`a3,q
lh�/vi��m����#:*п����"���H���p�ɍ��U��� P�$#U�FC� 2��6 �o&�"`��@#5(;Ŭߌ+%H;E�����/�lE�Ǣ�O*_ ����0��ͅ�z�[j@[�?vLW�-s3�z�r���.Ys*��T�����2�ݮK��R]�=={f���R�Rqםx�X~��l%{G�r�ݞ�5�Z��B'9��->�}�i��^&���qϝj�7�gp&;]
� S�-� b�&�eV+�v��3J�kq�DC�dl�g�S��U2Zb�MhR��S����u���7�V�}�+I�'l��rk�����=����mu��8Rߐ7�`��7���� ���D"��Cw���g��B����J���k�B�{&���죁��yeɝ��W�>���r���p��	�k�r���/�F4��`����녵��[xRƄ$n����.���!�/�w�.4�F�N���@{ML�nl,��mlps^���tq�Y�����z��]��yf�;n	�rd�7r�<mluw6�z�]t�t�gǭt��f��0?�?�yE��(3Fv���f�a�+᷊�+�)'%��h�~x4�3l.{�w2D���굙@m�ńZ����;����+X��t=y����1X%�
Jƥ�|��.2`|h
tӡ� #��
CK5ҿ�0*�R$
�%�p
a*�J&F����Q�8_����V \-�s��#<�<�b�ȑ�� gR,����ݞ�	�k҇�R7S�fyӷ))�g;�5�IJ<��3��l�X%{���O�5?/�R�,��#��j��{��̮�=9�����y�2�:�5ϧ�nu������	E�\)QbH��%H�|�f-J�)���O�[�4�K�E�W�L�����
���4���8��Oi�@�$\��Nt�˷~�E�W�J�4�EsS�4��2B�w�D�������`^�g=ƬDT%n�8��	�Y'3zQ���Y0��OW1��ʵ��r{�'����ӝ����
1r��	��X�A�<�;�>A�w���eh��{��{��B���ŃR"����2p{�1=T��9a�`�禰�"!Q)�*
W�"?���BD
�����R�����������ɩс�Q�,���0�OC	��7A(�C�$0!����զVB�V1C��
�.�Iȷ���B�����c᝸gp����	�¥�z�>��AFI�K�Q�)���0q"Y�bl�i�#��SW�J7@@���D�60VG��O�q�k�T�4�(��q*��=*���>G���H��I��؅���km�c�:�}ғn��5\���ܜ51�wn�fx�~�+�v�������~3貱��8rY�_��<EGN�$�R�&R�z�s�U�]�{�룹��^��C��nm<���}%��}J�MϚ!�}��ԡ�ϛ��ջ�i�sD�rƷ�Ŝ�\��L��\;G����f�<��,Υ.���|$�o��"u���!���Z��+N"}���k�-9�E�����Cv�k�k 7)����1�y[}[I[�l�6��u�:l���l-~_<����qGv�i����Zw�'m7�C�5ݹ�����/0@ͷ+��Ga0 �b��~��_�9@���
�,�j��7S�s���B������~��]?~��C
�[V����(�o����y��ŀ�r�Kk�O�}vQc�.���.�G�,e��b?E($ yR�o-���,�	dC���K�r�R����f�	�J?i�a_���s[�v�����y2_�07 \�Jf���k�������n�P�`G���՞kC��_���K��G��ٜ�0J��C�E�R_�3A�`����+�Vz3NU^��%�c���З���cȩ?#��)���m�.�R�#d��H�1��2T+�!9)|I5��P5�%�E4+Qk�jt�f5�	����f�+UkK� ���ۋ?��<0E��š9@!�BfЂIP��4�P�4�No"W���X<E�M�e�Op�ը�` �sv���e�U�{Ek��A��&Vh�k�d�Mt�#�P���"<�]�a�՛/X� X��	��TG`��.���%��E7�3ܿ}�$%����V�v�7D��7y7q&� ���!$k��PO0��D}�Nuǟ�m��@�T�b�h�q�c��>8:D�f�O~m�B�o�E&H\�A�1F�����3��1�A�K��i��HD��VI�9���{��;��q͕R?�|����Fhx����/'��)��_���K��ݞ�l�D���y��Zw4��-����	�t
�rA�'_�����Vb;�셽x��ٿȭ�%,{��Ҷu(-p�k�(]Y�vQQ�K�{3��JR�\�7p`-*ͅN~��q��i9�"���m�v	���@G�dm�9f-���<?ڹ�� فw��D66Z�����t�7�����Jȥ��D�ʙS�U�1?[���tL\���Cj��e�Ƞ®���B�kc��SRH���P�[%h���p�5����3c�Ϩ�r�f�sX��I�Q2��B��R�5Rf�
L��l��J�����'7W����h��`���N���'y�k'#37#�l�vH�n��>ႀ��a���Kɕ���9M�st��s))~��$�i�/��EY�	����h�37|�l[��4[`�4r]6/9�%�\~C���FV���O^�����u���`�`����]�[oc6��]��fG���3��F��p:�w�n���vw,�hb����{.�:�"y��(�iٯՌ%�{%�w"Q�8�I��]Ö�'�!&{���͗����&'x���[0����r�I���~^�E���<��[���"��L�RD)s��.���u<�^V��m���.��^�ɱE3�gjR>���ވ�t��N|P-0�1�eek/��|�g`�F���a�#������kc��-k]�d����O��-������Sc�{�s�[�����ں�;D�CE�Qܝt�C#)�k�9�)7Tr5s7ɳ	o��tuRA
ZK�ԇaJΖf�<��S�E���x��2�ֵ��n���Ç�ξ�����r�_Xv����)q�8(Sx���<���Kʠ��p���;<f�n}�tH�H�0_�#V���З�vĘhp��ܹi��d�z���{�J���Eec�5�:��L��d0����^9.r���%�#��E0��kH�׾�7S푊�W:M��? h8v�A��5yPf�|��N��w�W�m2]�go8S�=s�
�W>E{�gŴ����r0A��P'��Ր�M4-b�sB���f�M�����mKr�=��Rskm0�Z�巑��KWUU���=�TiP����*nO��;4��>_�����>8C���]���������������r����ma-�����P�����U2��Z�f�Jȫ�AA��7���r��`׸g�Y�P�6^w���RW�m�h��0ox�j��`��o�����"Ȱ�;��Y�#�33ţ��=]�����+�ìR�	�p+��Yt)�7N�	�p��
�z��:f���|� �}f�k�8+Ը����V1��upN"��J�%�n�Ĕ���e��	Y/�m	�A��dd�8B���$�|��2_�� 	7ـ ���S4�����C�&���[V��e� 
/�T[�0�����W�O�>}�Vy��X�������77㍕�qY�����Y�@�>_ۥ��@�t�����Ŀ.��5a|?{ �  Eɶ�C�i���>}Cm�&��Qp��ǆ{wqlEIx1������p^��6����BU;ԅ��`��4����W�~�V�y�n�1��TR8~��z}�������\}	y��f��+��գ
h.[-�U:4[���hE��AYf���t�"��qN��Qt������B���'$��e�!UYW�ow��c�f�D��ۺ�����SiX��(���-Ӑ�T�#�D���m7�H���,g���n��Q>�lM��]�p�X���iW}C^����a E%V�'p^z���˷%��2;��Ȩ�����<��i�J2N�VЄ�T5�~<�� ����11T�V]X�wF�c�D�)7�ꃑ�:��$Ry�H�a�����W�*V�8��H�	
���О��ء��n��+�U�1��Ю�}���|xv_L�Ƈ�t������	�M#T2�ؽ<��l����\�7�%5�Ϻ�?���˥�����.�����~�#������qi�︴�w\��;.m�[�N�!�w��;m�䖂z'��;
�#��N�;�Z���w�3��`���8���1�qi/︴w,r�;��}�{������_G�N�-�w��❜[�H�w�Q��ѥQ��K����"��\�  ��ϋ��~0������[~sƿA0��{5@u ��=�o�����؁�������ٚ@�H�@TE�w������@�l�0���o9�����������7������o&�����N�&�V����ud�#�k�_��z=+���L?�Y����������� ^֫S0�ʢ	p(��ڷ�,�(os�dA�>+܆?�o��
�8�k�9�4�i ��][$���pl���T���پ���) �I��� �E(���'���w��]������¿�����6���������m�Ϟ�p���~;g�ܲd��� �t#�=�T����	�PP�$ ����b+a�1�G�sD��rû�*�e�KT�o��w,�*0���k^��Q�� ?.fF�Z˿�7l�]���fm�I���=�J0� {�5`-�>pL?8: ̠K�O�~ͨa�~�88$��z`���ahP1�*SN@����ƀ�!���'�9���i4�>02|Nc��Ic�\3���n����߰ ��~�o�)P	�D��@��M�a�{��]��p.0�=��!!xj0 ��ă��?v���U�ΉR��s �7g���೼l�ew�m�4�5�|@K��gU!�~2�ďp!H�B���*���������O�Y�K�ޅ��h�d�x���x��Kp��iX6I���m��b/�dm��c��{c�_�o�::�������M'2;<���L�R���e���=�V�_�����g���]�l�^8`��/�\�]n����Nc�^r?y˙c�O�!�
i�8C�>��["��l��}u�?!j��C�r7��?32��//q#�6/K��M��[̈1\��]�\�k��^m��M~�`MÙ��c�I��:���0�:Ȋ�5=[��-�6��hX��m���n�Q˞��妑��'#�i5y�M��E���!��a������sq�.�٥Ɲ-,w��O��Ҭmz0�9���l�Y�0S��"��@2}NH>�u��[@���h*��Lմ��?K��Yw�|g	X��1
c�":TK�*��|1�*��Uh@�RD�FF)I�o���6Q�OM���n�9���,$��P�&�Q�����*�|z�.1&KD���q��?SP(źsEi���i�t.����QQ���:��U�	��9��ȱ���֖9Ȃ&ʶ���c݀��	�&1�9��^�
�4���j�.Z��DZ�Ҋ&+��&���I�!�w�J'�/P�}�\CkB
i�OS�9�G�H����YWo�]9Pz� vb�o���y����:�&Y}�G}���	j������Q���
�1��#�J�Ig<�+��� ���ƿ���XiG���Yuѯ��N?9�ԁ=c��$��:�g9sJE�����>�a��Z�{qr�����.�յ�z��h�Kpk.i��6��b7=&�c��ù�f��?Lg�R�k$1E�1�M�#@���q/�O�#{Zd�,G��^L9G4?�������[��	�T(��'|C	�Fj��_0Y�ٱ��7N�U��؉�n&aτ����~�ļK*��c�e#Y�h�X�'g�o�ǧ�`�:�M��R��t��<�ꕈӺo���\�(v�	�$ўZ K���자*�(z@v^�|\�dP�H�.	� <���t	�+�!��w�r�[6Z��+�W��`�������>�Ɏ��hŎa�W�N�3�b��,2�ùV�b�&A�?P�x���B)ΰ�#c���2!�n����Bե4�A��I9���難�sK����8×��5
D�x�~b@t��y���-ݐ3�S@h䠸S��H��a�A�')C��tW�1��y�I#�������G��������;�L����W9��ʣ(���d����[�ݺ
����V��f�m;v���@",�����d���6X���"�q�}x�+�V���ty��f��3��˂2l�D�l��qP�����}.�g�ed� �d�u�b8l|��2�M��S�lx�g��쓾��}���_/�:��S˜�&�50��:Bp��ýA7G������*�o�'<A��n$䩚�T�O$�H�������=���������ۈ�r*��W�;tt�T�Mx��N��, _��C/�zJ����� ���N��i��a+�[�����g��Y~��|y@����g��_���ϲ��� ��Y�߱���l��Z�W���>�eO~�˿�|��w/�׀���~մ�j��  �XA�_�S��XA��̨O���, ����y9�@a��_n���e������+��O���
���~���e������x���C^��]Mo;�YT~�H�D�̸8+�kwl��8�90sXl���M���$�!�����N���3��P�>yM�e��i1KIs��T��
���Y���܊�N����w�g�Ɖi=v��w9�����_3a�n�����/:���*��@���7%��D�ؒ��U�-�$=e�CjUz-���(:���c����l�l�Wy��U�w��/���j�X�E�3:����IM��_��S�"xP�y�Ԡ���(�m��S	�P~$ɫ���p�露���ñ��Pn��$�P�1�SR@� �x�5H�X噫E1��-��p�x��ꌕK��J�ʢj|^�!E;:�#
Vl�GDTS��ǔ�ٍ-7��Пe/����s���v���o᭗�?�Z0 %c�lP�WE92w.d�q��J�v����ab!�� P��o]�: �ӫ����_&}��E��''�
�H���E�7��w�Ey95���,�FO*4��O�ό�3��*��S���8`8��X��|�0�i��/�R���a����f�$��kb�
���&�tΘ�E�>�Ԁ� ���W�
G�&1�A?-�
�j� ��3�Sbbvo�―�i[�*��/a�Nzf�l�*�~`�!��R`��+��!UsM�"�@��qq��T/���<���@W���R�b�ǳ�S�[�m��v�)1��ֈi5s��U^Ң���N�;!�)Ȼ�K�Iq����J#1�Ď�����
�V��<� @����8��d�N��;d`5��cQ,9BԔB�XPld>��9�WRJ	V��i1��S�ыZ��D�H�����$���m;:�v�ul8j�p{PI��$�3��?��$P�5RJW����z����6�����"���$_�<˶az|�W���)�3*o�l��b"
���U��>+`���mO �D���1ءA��`��Eġ�}Ӯ9����#n5cz5TL}�'���h�'ɷ�Y�Y��C��N5Y?� k�� �4x�i�.�T��2G�/@-&NP�@��P�v�9qȥ�pU�t������S���KN"��X��к���Y1��bhi����-��U}N$W�g�S�����Z�R�Jl�37�/����e��q����L�Z�3��)뉼��I��9��O�4rˤuK�?d/V�D.~v���QJ|��H�J7v}ж�����_�6���5��,FLq�~%�p�q��ʀ�P�&O�'s�Ӊh���}�`�0���������©?��b��I�A�G| �i��!�U�#���� 3������y���`&p2Qx8p!�/�v� �3Ơ��=p�t����>�y�z(�������̜���؜2X��EF��rC���&��p��PfU�L�F��%��u� �5�mI��&�-3�L�4��&�>�<7]���sX�Tx�>�Scj9�5��x��xz�>���("�7LQ�V(R��̸PE�ճ�!�XNw5(@�+��(+E#��Z��'i������!I<�Aᆩ�����J^l�D-��G�k1g9��P ql#ضiZ�r�s{]b�n����V�9�Gt�*!s3���9��E�-^���Yʻs�{!�%�X�]tU�Y���5�����}��=��d�%��?�t���ת�S�Q`>�/gҒ��plŊ� s��[ׯf7�keq/r`��nwl�A����#O�K�Su���1��ǹ1��w�y ��2^��F��_�a#��<�����]f�]ly!��$�eNw	r�n�o�M�qKt��͵05�B6/S4냳��Zv{O��C��x���r��"[M�&�ڽ�hty~O�?8��)^�/�V��iֳ$8};��t���~��=]׋>�"[p���.�Vܬ��Q��ֳ1T�Pnf�X�>�ќI[k�Z{
!Z(4�zv���oۋ7��A?���N��D������� �G^A*�q�R�Cxe��
��G:[�~�'�:7���g�:��D�(�73���S����ZB��ɱ��9{{�c(�p5�AgX�v��fc�ʖƤO��O�H�Y�r����go|�=M��e[��D|<+>U�C��@}����I7���\��D��mlY����Ob���M����|���~�]���>s���aC �mc6���8D�#f�曚 �p}�����gC����6%�ѳ���u�G�'�B��V�N�^�3\��!�Pz?	wKE�afJ)!"���|��|)�=�i8ϒ�W	���O|�o���hx�R>�t���[a5��G�l��ح%�%���(!����&$�n0d�x$��0"@6餅l�XV!#�k�rqKȗ�)Se匰��v�O���G��Z�=Ҋ�	@n�z�v)��@�(�?C4r{��]ke?2O���w3z~(i2[��TȊ0�;�Eo��Z���bt����L����b�{�T��x)�f��|�T'���UC�#W�L<Oԑ�P�=40��
n
��I��,{�'�˹\��1��1^�-��}���8�-�L���V˵O��U3Τ����6���C�cy�~������V+H���r�j#f
�Q�XĚ����T xg��.��� �>z�2%���[6⩆Q�a�=��t@�-�J<�!7z|ЙM!�I�+q�"�|���VGV�)V�;�8>B��Q�c������k���o�[Iay��xod�*g���
��L��S��J\��i���N�xM�h&u�ց�K���R�ѡM��Q��4��Ù�,�F���c�D ��A�^�eߴ�8"�NH���cC\��E*m����p�1��n��B��1���wz���\��r�{.��I��R�`��E�1�j?'��,!!��a�n�h�}�0���#>��:U����"�g��a�R0U_i75�L`n�FN{8P�����<H�@JW�$���O�������SN�AJ� ���M��^=��w���h����k�J�H��+�q�w�&]�q��lX��lR�r!$6��:�)����ö͕v(�M���>�/�Z;]ޘg��tP��jT����j�,�+��`'����C�y�C,=����.�mbBNr�V�����}�+yx���f��D�(��ʮ�O����M�����gS�'k_��CM�G�}�mNH�k��lCF���"����=kI��:�7�滢���}����◤����⋑�5�>��F��>T��Wm�C7x2}�ZP�\(5�u����n"~�r��?��q췸r����o���z��k�
�i.@��w-+�Ͼ#Vp��W����)߽qb��L{pPmBm�Nǧ���_��S~h�~���}����Id��X�
���9bf�˾jhd=)�BP�3+g�eK�L��q7/���,��ܟ-��/߳}�M_Q���v<o�ϊu��,MJ������4��&�Äs@T�]r��(si�!Kg;�,G�G��˂���Z j��.���Rۮ���Lt׌V��L<�H$ď��՘�"�
�*�J�b�×����~�q��,�]��k9�=�����d7�z~�ȁ�b��w^�#5�l��Ҧ��Ƃ�����R�΍j|k�G+ۤ��@[aX�z%r��1Y�M�:rF�S��R�DI�+�������դ�E}��o��A��L�vM�����%�j	�t�����g�b� �P����VۢV��ɔ�c��='��o�ߜa]W?RN����H_0e���3@�����*���O	.�G��a���Q&D��LS?�
�l2�r,+7��+�L9�0�D������f�(uZb~SZC@K�Ú����)`:i��ܯSPR9P��T�tF$��<L`z�l\>��'F5����b��Z��F����cy4�δ�)��$C*������W֓:t#��� fD���g^4����!2���·oa_e�-M��	=
��	���O��lmF�|��y-⬶^p�7�#dD5v$ϗ�!�7��ל���J����3�,z�U�nKV��f��֚��٤"���%3�G7s���gs�C���blo��Xɔw'�&��-�gR�_X[�FQϜ��tLo�.�<�)ϣ���V0p��}=�z�4�%ǜ�A2���3x4,��f`����ҜI�,�C���oȷ&ٸX:D�M��3����iV�V�M����#H��4�O�V��"L3��!�1&cu^c$j�|36ڄ��s��iDq���>�����#޶�2�-�FT�q���R�p� 	^������� ����y�?�Ȣ.�LI�',69���J��[��B�ANz?��8�k�^��w��[�V��x��a��{�@����B�<7��r�	N�1�:�<�/%O��܋k4��:mJ�� ���ĳ���7V6�=xi�ɂ�/�u}Q*Gn�ġ��� �}h�R��so���؊u9b3�Hx҇@�T��kRuI������ �7�8w��_;c���,���}+E��g/�GI'�HM:1�XL����؋�+�����V���6ϛ�HGy��,wQ��ܝ�a���y).�n@|�6p�VL�Sf<1 ݊I�B��>�Up�u�~/��N}$��f�*:�d}"b��XG:ޤ>;��f���]
��j�kb���p�Y�k�̠�Q�`��u��N�����	�a�q�}�QS?N�ƞ��t��[��q�9���iN�j�M������Y5���f�����G��&�{�.B��z;����x�a&�󅣛��Q��6�I�����[�����I��+m�����F��?YR�B��+��9CMQ���i�A9�w��Q9��0�Tz�;%6@<��z\�8�0	}��e��m�H�ְ�:�k�	��$�+�
���?�}��e��g���d"����s���7����F�c'o	}�m����>�����5"�/壆�����������M���_���Vx�̝P+�]]�M˙ʓ�5Z��e!1 >Ǝ�!�<��\ ?��6ekW-]�q ������\	n�ۉA�xVŪiB�Ê�Fb��bn����W�F�����2�~0���{���j	�fo�K�ݫ����РƩ���/m]բ��G��=��qFZC:s�����:��_P�L����&�{����%����|Cֺ���y��}�yf���5W���!�1h. �u���/�N�Ci�U=YO��y�[���J�6'5Ӓ�q5�j�	Q42?��>�(W�L����g��^&�)u
�N8^�Bx��)�"?�Z��g�=���oJ��B�mF=X���O�ԅ����qn���NBV���	�[�3[�~.�i^�W�5����d=�k#%S��1�7��ܗb��\��j���iMs�C�F��R�j�@L�~ۣ�s��-�L�'���%�����בַ����;�5�cz���6wM6ޞ�%���9J�i��+
�h�IR�l�P���lg&�xRl�P�Ȕ�`�25/���6�e�K���:#	2�fM �/\RlM���%�Z���V�36Oä�kv�%������䌧7g��,Seb�}SJ�db=m���_�E�N#H���r}� �����w���񵞮�U+V��"+�<�V����eG���i�t�yc���Ii[I3�8��y��oL#�E�:95;�>G���S�<�'�W���+1.2��F�r�&����7�3S��E��>\�S�|����D�"[���$M82��3�(��[�V�1�9��� G���7D �CK�	8U���1c6ې���TK
�Tf�)�Y[ƈ��M2OE�L'2�L�	�뤈I(;������{o����s��?�y��l���Z������w�k�}�曯�3�+���0�.S��h��6�IxA�N��I�s��-K!��e�-m��4�R��4���iKE��@�.�,��%5��ϵ�O��C��Tk�nk=}jV�f�v��Bsu��C}�B�B�Ǥjr����.�ٚ�Is�S��G�?�����$a<ڮ_��t�h�zp��!B/�OA|�~�ݵ�{r�<>��$B���-ai?�֘�.���̱����7�f1��5�X�O���r�%��l�����5|8%�*0�ms��CVvV��Q|�� }C�݁g�Ǖ���:�K�N�)�g�.���L���V�5�v�	ͩyt�%����6K�Ԡ��1�ؒ�IaB.�U,��P����rݺ �̌N���^��p�u �T�q��G��p��Ĥ�"�+8?ᤋ`�1񭅅1\2�{Y$���@W���Rߔ4��ʇ>f��5YC�P�mxt+�E������S& ����q��H�̺(��)��2�:ɹ���=���l���2l�Q���6�i(1�?��n���;�&]��[-��ϲ|p^/��
��-�<l���J�L/e�k��J�o$��D���ǚ_���h���%^�vOìթ�Ya�v����_C���]D�^W|��e��G�1�1�����_��������n`/�*�Į����~�`�t��E=�;7E�c�T2�ҙ�4`7_r3����5�3��ɦ	)���������>��,����}���F�t�!a$�N��d@�c��~[��q�W�g��m�����'���2��7L��-���&f�秝}��뛪��xj�:�h�>���rJ)���|<S��i����.�D��;'��Z��-�g��]6�7��L�K��f�Q�V���V쓪���Z�ڙ���7�3�����\نsӯy^��k�m���wg�U��Mj��ܼZ��="���g�{���֝7�!��9�B�@mc��QN)�b��|�^�	��ٷ�x���m����
ˏ�\�(7o�K�m��u?U����{5:�'ÍG��6�����Ò�e&m�z�����8EF�yh|��ĕ����/._��q�1�ǹ��f8�]�o�m��]Ye�W�ː�ȥI�Gc]��L�!�Z�,�u�d��FV2�l�����?0��4�ev��i�����f/����|�XG�m��?��I#�*���9��J���h�x��V2�4|�K�˗���T�.I#_,!m�:9Uhϊ4|�H��U�q�*�dȷP}�'�?����%�Ѳ ��nFj:S����_��u/�"��=?�a�y���}W��]e�����.��������L���VO��L�����lQsz�U�;ɉ?2�;�~��9���@��8�<�GL�'z����]��-_���X��ᵝt�n�x9�d�� �)���R���h�3ݬ����?`�]h�3������|���3��v��.��߻��R�_b�������� 	��{.�c�w|D��3\O��3�4�$W5t__��𚠹��86�k�^3����ýE�jpߚ��BD����r�������2Nd���I'�mM��K���X��z���&�H���\qs�1��{-�*Q��s�/?ҧ���&���9��^�5��]�|���1�nyMO�5��^���#��2	[Uk��tuq��y׈葮jy9�ӵ{��p�d�6�!XnD��lV.1�)/��E9��>&���������\~	C�;r�%����ǥq����*>^$�>�5��u@g������|�+����g�����!��os�n����n;/^Kަ��5�r����K�_���M<o�T���<�m� 0h]EL���b�u�X|s���\�3�H����XV���{�<q��5+S���s)9�t7gH'5��t��;���wK#��ޞ��ǟ���:9��f���KW}����	���JP�a�c�����]�.�Χj{7_�['b)h۲�����"e�����������-�ցf>�zr�)'�u
��m���u7��	�M~ϯQ��$�WZiFm����O����C�m�9o�e�N��^t ��f���+��LG�:��RuX����7=���̫{J��9���3��w����_x������sHBi��&��Ϸ+\;BLY���Տw�/h��6�		6)�䈐��s���To�]e��JA:)r�/Y�`q�l?F��n�3��l���y�M�#^��F�q̚}�Đa�n����饽�����%�}�D]�������/1�W��xwlޠ���-ݕ�!�g�G7�ڣȑ��y�R��������6E�"��`�������-���[��X�
1P#7��'��mq��X�/$I�X��zN���_2z�d�a���K�3�o&4�^y�8���L�B��˶s��[8M��]�CB7���i&M*lx��*����`�q��!z��\�M��!��7���������TWG�$�ͯ?��S��Θ[����lA�o�c���[w�MsMZf��Է�?�.O�O���#���N��9g�>NvÏ����:6�6��Ǚ�p���W�18=a,+�7z�A���zҐѶ�sУnѳ��S�gߤo`���j�wS'H��-y���ӿ�<;��4�Y'OBp@Fli�ҩV�A��
�=y9�kq��4��ROY:6���nO��`a�[���V+���~L���oيj��CxG��Ζ� ���eQ�jJ�l�DHJ�,cxX�#Ly���AUl[��WB%,�j	/M��.|��7!f�=}7|�C�"��A�^��ث�����&��TI���K��L��Ud��z)�K��{醅��h������=b��qSs�]tve`�g���"�P���~��8�|�μ��>�r��Ի�'��M�tD��e����H412 4G��XJ1�;��m��i�� xţrmC}�\UZy�������!��Vg��%�,��E�7�z޾/��ZV�j�cgXsᾁ̘�^#����Ro$DJ���i�ؐՔ�_�8����Z���ԔW��+z�ͬ��o�xD,@�%�!՟��@s�Mi���I6�[��o<�vn�u�,׳�U���Caa�nm��T�ŧ;lz�bP��ѯ��.��\.Y�Os����6*�}�}g��4���t��]��d��������q���ӗ�X.�-��˥�2�l�\�,���<1�r�w�>ю��?8e�e.���d�r�m�.���7��<U��%MqY�q����I�k�͞��rɫ�)V�S�^����0��y��C���W��z(C�{2 �ҩ�n�򞴉O���]�d��1ɦFԤ��7�Z���Z�e�������ϯ]�v��i###AAA�B���GF`�I�Vl#�@$�v$�	BH$�"$ m��0BHB@Qea���  &�JA��U �[ &�0� �!Z� "�C �?���$La����B0H�AT;�)@0@�ю  S�U�U�t�zBE���� f
VG�`��ݢ5	"�	�E�@7�$!@�F�B�� � `n�܄�F�Z`^�LB��J�Z����Q٨hT��ی��$� ̅�}h�hI �z5��H@ �Ա���<��s+��Yhk� �~�B��)`���a�1� 68���� �X��D�C�Ek�s�Q��
PG��@�8@�)@�@�@���P���T j �%5%;���������������/""�~���7ZZZkkk���"�Ȉ�� �
S�w��SS��)������.��d����r|#߃4���D�;�����d�+@F"����8 %Y����lAg�i�i3�cmYP�I���Ix�P Ï�Ư)��?��T�Q�����o95~���Y����]�߿��~��@F$���	3K8n���E^���=GW�����	d���dU�"�}�م ���.n�(F�#�_����$V�Y��rm =lNvߴ��)u�Ƴib$�	1�C��|��#��������M�wY\���]�н��谗�%�|��!�ny�Ò��`^�6A�ʰ�;$쭂d��0||n*�_|J���Ԉ&�p�_�u����L�5ޏ[�%��<3N��;̙n^��5Zs3�N�"4�0����u�=����:Z�Nh���u!�i�Q���=W�T{��7ܝ�:���+n�;i"�=VmAp�ɂ�O��а��g-�1Yz�ȓ���Ҭ�B�D;q��)������t�*����y��J����w+�H~��m�3	a��g&(▬�Ի�WR���E�wo�۾A���ن-3���>��-��Jѽ5�;�B����(���n����֙�x7]QZ%���H�����/��*9�Ez��ݠ���b��P.��yK��9�����ʎ��"2���{x�7�~jRs�1"84s�U�-��#�iq��ž=@��L�x�\�P����z{�AW��9�Ɏ��k9.������ �cI,ffffff�-�X3�e133333���,��}��g��<������^��#;��Ȣ��ʯ;�R�{���6�_�g�"z�zm'�UD�sM��O�0��jc�kd�,�\>;�"ĺ,*�#�[F5H�hJ�P����f�����[	�o_�q�(p$�"��Dm�.���"�'���&S��tޓ��:��6�`�P�G�둜��#�?�߱��t��N������6x��\P������2B)��5 9�y!B��#�M����Yg�ky�lG��&3�Q�M2�pE	�v�́/ܷ<�5�3%���rB+tb,�d�PB2tk=��&v�Vj��Q<J�~����x�T*��M�|j�"`�0�*��uE�r` �sW�`!�Q�&\���O��}P������߷H1�7:��o��6y���\9��o"X�[�D˸�V�N�SVWQ:u�Т���5������Td��[�iX����.����2�ȑal�){����۟���P����,�Q��H'*v�b�7:L> dޗ��w���ۿ�U���4�cb���������N����ʧ;�\i�i��yf��J&Y�#�Z�^b����0{�ˤ�$����]��Of ȍ9���`Jp�e:t�f�����ֲ�y�@>�;>�3d�K�ZP��c�����F+\����p9а%�jB��!�-;�җ��#j��L�e�l�Zx�m6�b��I��EE��m2Z5r�B٤�
r�ڥ��:��I	9W�!�q��-y'���S9�}�`C8�����U*Ȁm@�(��Iq�-Y�`��@�u�feeb�ꦊx	�n�T��ޒ�tZTzz-�i�Di�М�<�-,E�W�0Z�'��Q��ݰ�W�a �N� L:=�q� �x��R��ҧ��`fC�Ep��7"G�+�>�f)�&T9)TΈ2�E��BJ�����34ݩ����#1TM��:�TX<yUn�Eo���Z�m񮀬�V�зe2�߳"���$������fK�"�My&_jM����ߵ8�|e���T��!e(ӱ�9? ���@�}X1S�J��\#��,����� �,mfu�7X���삑�7V��*O��1��¥��Vq�W7T���N�?G}SiC�cGl��ʾFc6U[���^�@'ta�A�@�(��pƶ�������������V�Qd�ŝ,���;$�$:�Rs>�����v�B���A�m�oyz]sh��FM��u�0f ���YU����=�a �n>���6u�{�(I�Y��V�MS�/H0�\4��O>�<NW�f���ɒ�,��Х�W���BtֽD��M�%�9����<�f*x�Qi��v�y���˻e�th}�ۿW<~�O){��t5[.��+Q3nzvX�.-��gw�F�����7���c��?Rcʆ'�W�SE�Y��;��y1��3z�G˕��}!����ӨB�p��� �y}kSkI{Eޭ�cs#���sK�ӗ�m�t�W���	���}�	�ڙ���ƌ��y�����Ԗ��l���tI�+��^S�w�c����'��U,��\Pw�a��)#�,{A�lX�h�t(�L�3Q�|��F>�1P�s��Om=�X�{#H��ȨtI��*=����.5�V2>�̚7�,�++#��zז���Z���TkdOe��.��Z|��e
�Io���C�'�░�^'Ӫ�N��.�e�B)�f,1�s����VO�BK�#�T�e�	��0cd�:��%�ų,�Εd�i�j��dK�\V��^">o�+���p=G�-��e��-�Բ{��l� ��W{;W+Q#�#�=����=�:����^��sތuIEP]�Z54%��{�@Đ9u*Z;���UL+������;6�`&��f�Ibv9i�	t���i�K�g8�ƪ�yV��3i|���Ϊ��͇�X��[���e��J�~&��E��~K =�!��"lFa����9d��>9/Mv��'#���_hMS�Es�E��G{4M���[�	J?[��L�����t�D�Ù��������g�´39�z�G�TF�����36NX*���i��y����uŗx<��9��|.(�"�ٳ%�B.w4�,-�|���*�җpoD��~H*`@J���O�N��+*b�ƕ���#1�6l�`��w=g*�a�&�R6�jv�΢p%7�)�e|0�\y�l���>*?��0u�7��a�֭�D(�Ed{�����Io��AY-�Po2�6���:c���$*��Yl|�9e,j��*rXP���ﻋ���hR�%�y�	��^)kj)��=��_�ى����߀π�j����ʀ[��
�a�e�� �#��睕�i�W�^��Ī]��������|	�X�����������-2�"���F5�\D��r�׌�G�X��6����������A��J�`�f��kv�=d��>�l������Pne��\`x��
EG�g"K��;ɽ�;�ql�^���р��;�Z�e���3�Q�u��a�ڞ]�h����oN�K�D����,��~�>m�WFw���텞�%Il��D
_�.�f"Ty]D��;
=G\䤣�tZ
�#Ya�g	S�s�,�_V��(����Ꜿ�����2!8�q��k���6�Q���y�1���Y�\���������㱆��cPҍ�4:�yT�$��]���M�{�M��	Ү����a5ތ-a*Ԗ-�p/id��i����1�N���C-����u0����]7~D�H��'1��p���Ӫ�e�Q�UtR:r���J[9��3�<2�;>��m�櫉��8pR]�;啶���'DsV"-���>��d����x2�.2P��"��56�Fl?�&�$�诰�Q2����#W�8���@.��lFj��k�1Âv�O@)��HW��>���7',��"�ՌY�� f�����!�Z��n���Wz�as�O��m�dgذ`�/���޽���������Х�d�>�䎉x�N[�d���I�;�:z���{C�C0AJ�d�v�7��2}�hɟw�"5�D�i���06�<�nCd���Br�L���v<6�p4o��9���Fg[�S$x�՟�n�Qv�C�CF�"9��a��(x�w�����3�5L�.~�ڕ�&�w���u�]�ysf5_ʕ|jz^�L�lR�O��d���D�k�n�hfX�$�����c��3�լ�68׳+t����+��Im����O߬Ǵ�����Ǵ�=�G����HA0�A��ҏW�4\^n��:7�D����>�j�=70g>���Dh����$�>�L��ѽg�xP
�zC?``#�?Sī��������������|7�:�g8y�N��~�������꾡�}Sظ�}�/�!��������Y�k��� @��_���b��G����Z�����-����2꿴e��  �\��5\m�0��k$��uS���ԌW4�w�� u'����8sh���n�YB�*������MK��-�#��e#�5�ӅLXA��Ex������EX��>C��)?;@�|ʠ�����	`�_y$�k11���R_=M��j��j��P�����m��\&�K��F	Ǵ&"�]g���q� �dg(m��K�4�E:�(/$r��㻰)!Tr�a0 ����ϰ@�h@3� լ�HE��(_Щ aŅ��YS�f����4��Ⱥ�������Nk-V����WJ9�jx7r�be,�AJ(?�t���c�0˂=̀0�4R��~��y�0e���OI=��v���^�
-�ɠ��U�͆?��8��2JC9Vn��"�Q���"���%|p�~�^�`�P�C���D����RjS�,.�RA?#D���/E�P�;@i��H�#�t!E�<�/�"_p�,bQ>/D̡%fR�K'�B��$z�U�i��A-$n���F�,t:����@�!�'�k��/f�0���/�~s����6`�c��e� �(�̜�KD�	����NӃ2`�E���w^i<�h���)��0
�Sa�KN�_��x�)�C��D��pş>��l����T[}=��ʕx$}�0��R�MD%�:0L?eB��-	hG �Y'ۙ֊�9�$�%MI�oż<K,��=���x�������m���-�{��v��VJf����/Vv=��S�+��4�bY<i���~�;G�y2WI� -�'Ĩ�Ĥ�G����� -]"�|��j����� )�3!W�2�c�����mf��8�>��Ž�1�y�<F�,!#W79�}.T��԰�T�(t$�0������Qe�Yzp�Z"Y�E����:_�b�Bŀ$�y�8�a�4Lj�L
�I��qy�9��i�J�܆�U-j�^�ȹ��-73������Y�)��NM�P��Y�-SjL�5�]���D��D�z��ޑ�6�~l����X����1�K��]��v�Ⱦ�� s���]�0�J��x��X��5Z���<��W�ػ��_S��{"y<YG�w$��U�J���v���dm��ڌ�*sz����vf� ����.�.y��)���I�u�t��,�����jr�u�I��n^�>%��pQ�����yZ�s�B���[O$�Ã��kC����t~\0�Gc�Ecq����|tk���P_R;S�W��[
�FC�������Ap�V�J��r��}6�^�!F+13$�ImI��Ju��ZF�b���9*�1�k�+��`>L��o�?���ѴE�e��.˙⊶�ɴwdT,Ի��.^���=f�}3n�7ܺ-#��%�g���I�av�df����@/�!���$�#uԸ��o(�}�|Ţ�.u������B�jhK ��LB��9���Z�7�%C�5�g�Cի�m�G+�����q�r�O�H�IHz|�������őM�Ť �(3z���C���s���k�B 	Q?J�$^�e���ƴ��g���6tL�w�J�K?,��%~��ؼ]-i�-H�����N��~|�}t��C��9Z�E�;9-7�H�y�(�+މ#�^&E�Y	��n���^a�I��z���W��e����B�{ӡ�O���ؗ;��ӗ�ǿ8'wC�ZJ��"^��F�?o�*�O�w�u�_����d�����E|���:�RDl�����x���nl��6e"k�Mmgwp8 �^��[��H��(F���V �`n�~r����/l/S�F�[�^R���l�u�mgqpgхN�'��I[�h��»���۟{���7%-�?<|u�b�XSi-�-z}-���2X:�~� m�Ŷ�l��˹�F�\+����,��d�T?�u��1�%��Q���ӮUr��5Q��BgF;Q�G�K���\%�n���zאݕ=
K�M
�Z�Nr����T������oN�� WU��i��{<j#�Ѳ�t~G�:���D$bue��x����L<���n�
�|n�z���:��#��,n4@��U����Ji?��,�o�C�ѾR�[�JV�C�)�Sd�߅f�t�O(5���C���� Ⱦ
qϧ.>�dl���.n7۔u��L;��0t��m:P,�v�Y�8h�'(Th�G�V���.<�Q���q��߁����4�üJ ~n�Q~�Tί�X� 皰.�Ғ�Mut�=T���K��PcE4 e澴�*40#�TX*|TѾ����(�P9�&N���uP(�L�K��啕�;��&uxQ���O#t�bѴ���kvS0;�lt�U�P���_��\p�E�k�M1�Ϯ�\�f��Jj���M����AHG3�~�|cy0�F�+��Uk@��^	j�f��z��F������F|������DBJ�Ű�V�yF�ܱ�<:;�8Z�������H-�S�ZM;k�&y�$\R8�֟�8�^�9)y;'EK�}��Ǝ�	vb��8��f��4��Rs�L]���>6�S�A��j v����2$�=K�Ii�	e�s���O�@L�[�5{�<��I��i���r�B��8��D:�ܫt_�S)�y`�'�9+���;�$�����%�#�cO�:�kD�H��/d����O6qI�3}���'��d��y/	w����Ȣ���(�ޏ*�t}2Ɓ� [��>U�x��n�y^}2��|S���`��9�&�]y2�&��8OR���x���g೜���X.O:2��Vm���>;.RI��ލB�-;�=-uM=μ;X�Okl'�ı�	T�hU���O�sq�~{	3T��_Ҟ�A(�B��o��/�_0�	�vQ�Z[h)!�i�gu�`Rl2>B��B$BIxm9s��]�=0*F�N<v�K�CB����׉	z�{�������k�F
��:���a�6�  �N?������E��B�^RZ���&�,�m@�(�u�`M�|6)�u��^ $�ɊX	ē�����d��7Y�֥�p�/a�2|�B� �o�:9�vL���]�����|�(��s$aBD��'#_��O���M(:a�}�Ovc�8!4���"凧L(�!���z3\U� ��+l�B�٥��`��`�b��	�E�,�o%m�<&UA��nR@tS����E�淼m����]cHQb����|���<���;�g����1��8�2�����U�B�)����zv�:B���*�${��B5R^���l��������aƝ��7��i�hhm��O�/i:�u��I�OS6t<�}� z�.zn`	��dޣ
M������ԃ�!�'(�4&����H�w74�[A�Ϊ�L��D<7�@�,:|"k@�\��!�g�q�/��AG���	�)����ޟ�֑���6�(�~�jדTF���(�߮�/�9c�RM�?��bt�Ū^�\��ݦ�al���1�:b�#�������``>�tc��ρ�Z�ׂN���5�tG5ޤW6`���6�j��M�R�؋y����v���7LV�	���J��z��.~�~�[���4Z�C�p��3�B��QIa�����RD+QjI���Nאo)�I���w�p��9$B�q�/� }���z��j@i���V��?�o��N?���O_L��vͿ6 ��X�4l�~6��a�����?6Q0l��`�4�����a������(��P�?60lD�6����r��a��֟�Ȱ?6�Y6l ��l�@��ٰ����y���/���1�_�~a�@��"���W��/�Z��_�)�˟c����@�g�������φ�����c�6^oX�^l�?Ǩ~a�P9�"����1�_|��e��u�����6�a�g��/�?�;�Џ�������U�@��������_�!������C�{��o������c�~�)��b߈���>ͷ���4_���}����(k�/�2y��'�G��}}�+נD#����?�o0�����D���gDdB~|������X2�ñ5c&���h�o'YJ�5�,ss���Z�ľ����������~Xq;kG�?t��\>��\/�?������������%̀AOUA��{B�����! A�b0`�O3 (��H$b������hB�? |�ג�>s�?�8@S��Ⱦ!����c�u>�p̌U+��s5�{@U��!�ڟ�P�u�Y�����@`( ��a�7�  H�D��R�]�s��uAP���G�!ֵ*�>�X�(;4F�p[��
x#����s[��.���!t�>�@X;�%Lҭ�34��,�� r�s4bYl�Y�e��.�c4`ZƂ�G�˓Y��hC���.��� QXY(���ϠN0:=�� i� U�2V`���8���q����?���4r�~>~9�(�(������5�ʜ�Q��������qD'��hYUM�HYU���R����W���!ta�1��୤�o|��H̤|��́���^ۗک-�7Vړ]���_Sׄ��yZ�0fI/O�ˏ�?�'��^��[����(�y[�,g�u��U���9_�Λ����,�Z�"���R���$%ji����<h���l;
�VU���aŹo���[��x��A�(E��[*H������J1�Iy#ئ��A�$�IS۰{�R��d�s�^� \��)�."�p��]3g�48�(��K��WM���ڴ�sa�d�+��W���fF��6��'�'�q��q?I��p�y�����H�3VG�UB�S	�)ڥ�1������+������Q�t5�L����2m̗��J�U�S�ᖛi#��֕S����g7�tG$	Ċ֪8�%�����etT�T^O�e�WK��m/ʂz��$?��T��+��.�C`1�t�>����[��Y��6�v[�Ǚ���21�h��Y�'�̄�s�S�6a�0aD�;hq!ť���r?Dn�z;-e���t{����B͉���i�eD��M;���F�q��!M\Z�{��|9���z�~��c�"y�S:RT�"T�'�8Nه�w�hU���L����hC׌�џF���
Sa1�%]�X��68�	�	wgFEX%#����@'8�T�IhI/9W�
ہ��ezj0��n��JZX3ӆ�`A>������ I���a���Ǵ�90N�;�T�B4A6G�.�=6ix�KyT&+���(vM�Ϗ sA6]�HD7�}f�-P��D�>�D��j'��R����l���e��(L���r�6�ݡF���\P��"uN�3\L�Q��f��+רj3l�����.4�7����%�̴��U��<M���Ҕ�V�"��W 8޽Zw�7���̜�`zb��NjO��������{�t��\�D��:3H/�Kk�g�B.̮||?���.�Z:Hs�\Ş��0,�JXԋ�<�4^���b4���n�DG;ԩ�I)Dٸ��]�/���@P]\�!~@a������M���_�M���wC����\��8�`���0u]��Iu&���x�ͣ�,�`�$AW���,Q�J@Զ�:��_�5��߃�t����E�Ow�I�:N��?�й��1@{���BM�� �{�<S� �!�����������X��Z���sk�@^,��_ 3�,5`d�(���%V+�O2����?���u8-}W��0(B*=��1-e�|��ؐΰ�k��`-�]J�1��6u�{�29�����è��G�|��n��%�U/�z<T���1�p#�vq-}�|�!�St���֠��Wt�Z�3�f�oٺR�__01_�cNu�^���vUS��ԟ��L�!o|��0�uIܴ���K~�Q�w�]��7Ά4�v��H>�KK��
�^�㨨��L�C�"T�� v��U���i�y?�Ş���m�ƕ�8�U3f�g��-B���L,��+��c���n����mWJ��/@��an֮��S�xY�\��|�{dscڲ��j�;�V�rGm��a��=�Ugg7g��oWKW���nt��c!����8�%k�G�Ϗ��}����<���<��`����{���R���m����~�A��?���u7���~~�o'貟����̋~��?�ȟƐ�O��gn�3G�ٟ��3W�i�l�������i��=�����?���=t��1�������G���kh�&˳��6O�M�������N����w;�k{��=��.�m����~￿�����o{�[��������  �\����m��0��Ǯ��풑�����J���^E����d��B���&P8��������B0JAS�XC��1/"��P�[�g����������[������G�s� �7�Asu�`}�z3�-��S����-u2t��.�MH�ܔ-<���H������R�on��|2%������x{w~F�+;sv� V?�ۻW8�����і��}\�!���V��ک��ة���*Y����b*����\�3�l6��OL�)09��k��@|�������9����y��ibƈ#"i���a�#�����j�|"�~u9�M�?�!��y����
�1�8�Ī�C��Q�Ex�����7��>9�Bd��ڞ�=c
�q4�l9H�&p:�zZ���4r ���C2���6)�A˽	u����h�+�j쀰5d��Of���_f��µH��&�z�>7O�T��@����2GH����xU��] �!Ǘ҅i��E�:�K����!n�x���_ߗ�RN����XG~���M��iPbOhf	xt�����iº��.]mg�x^�6����e9�fiA�P��b ���VR��A��	+T�5�Amg܋�Ü��+v:p���g�&FdE��ao�x�G�iO+Qo�i�^"s��F���k��'�w�\q��]&qy���XX���&�������ƽ�a��z��[ƜGl���N4���J�v��S�����[z�A��7Rtf?pr9rq�J�Ђ�n��Z�Ilu�e[j_�ϟ���/�*�A)~uPݗ����z�F/�Uw���c#��W-|�Ya[�x<�������D/��禋�S�3�i\���C�p�i:�́^m��C.�$�[pό�.��w.��*�tB�;��	���M9��j��=n���䠤CY�\o�%�V]�Jz w�7�=�+S�g��B�%�|"W�mo�*��8q9ḥ@�ɏ|��s�"��Xf��`�z�,uL�YVI��g.��<]Pd)e{L�x`����u}7z̊Z`����1������-���s�AK*�9; ���|U.���o�$S*����y��w�ۖ��5rC6��8Ԝ�%�V)rNHu���Tڙe���Ռ���c��^�l(�������?�m�����Z6a��5�Z�?)?w�w�ғn��\F'�"S�?��h��`���>|�g8�!}�����p����N�֍��3޶&+�*�-SM�7+Jwu���C��)Ŷ�谇���A��4�[H�S��Tx}/������9�uE�)�\�(g�-�#0b�p�+9�r�,�Ջ�e��x?�3��L�P(��e�2���a�qҠ�=���� �Q� ��6��X�+��aFw����'�Z��M�NP���4�p�Ԕ�z��-Os2��M�g*���C��Z+r�R�#R���~}��`R��?#0#�#~��Q�X��Q��`'d��BH����͎Z�.�9���	�Hç�,��젋�vK\�M�D��W�o"�C�p6J����)҇@�;,����҃G��	gd�GB���T�I'Q�_j��d6)��������P ��C`?}T��hfw�yG�SԏY x6{��@Z=��� �B�c�<��iuX�O���ǀ�.!X�	 &����(�1\�GE< �)�>e�3�-j��z\ʠ)�|�;�l%@�Y�Y��$#� 2p��)E���:������ �;�#{ښ{%��T��T��gp�6t��V�C�{Ha��nwtA�j�0K�^d��k���wHkj�����u���-^��qf����D�W*���&���B!gv�������X
��Iu�+�'m�uÄ!?N�Hqh�r�6+�a�� 9`.7�r�Ӊg<>���(z�%�Y�z[�є슅f����^9d�"x�#�P�@�)䷎7��{�E�날��=���M`��l"��l2	��|Eoܮl���~�ͳu��+1Pv �=?���O
%Qu�Y�C �({6a�NԈ �D6��nM_`�����=@��~�h�-]�J�7��햢�j�Ȇ���$�(Dw������>&o����$�o	(�נy܆Sb�J²���cԧ�7#H��{�㇁��\�{�Y����J)�޲����Ȋm0���G2�\����&�)��TAO�ҮM&Rsuޕ�Ҧr��I������[�w�Vd����э7�V�����e���ًS=�����p���䥤�,�_��e��k�Q]��~������ݚ�%�>�k�y�<!�[;�`��:V5��g�B�;=�����I0��npڜd�X��&�p4�͙sv�Q�V�T� (y&r���8>�Z%��`�X����u�q�!�Z�I�B:r�����{�(iz�E�����9��a͗衳��2�U��ډ�����k��'38��D/N�k7�5
�D�+��
m��"Q�+�_6�U���hu�A���U�ŋE�/�S�T<X(
�J��)F�H6�Qj�.�B�ާ��nMjc[CikB�M�*%�\�o;��&tp�I�}�|YB�o6nV]�N5��:u�d�/Q^RQUN�3W)2�������`N�y��	�j��q��7KT�pe9`����B� o̘ ���/K��	�Z=PDf���]�-Pz]��5�+�P��{D��a���������,�$6%�\��w�R�q�{Yqԭ�o���v�$�㋳����ȵf�����;\��b��rȣ_9Ƥ>pS�{��o9T�2)���!��2[���z��4��(��%պ��hpՓ߫p�Υ��J�N����;T�ٱ˖5�7�PK=����f�A3�� /^�ᰨm�)�
��6D �������_��!ZGcR������^ys]��3�Ԇ_��7���;��	k5ۧ���Q��@���͂_��t��YU*5�bXΆ���ZdW;����i&Ռ*���� S|�L �CK�tI�`�333�%Y��bf��,fYd133333X���kW�gjڮ���ݝ�s�|��K���<��q��lvdښV��M��U]:����X^W��p30[5�<fD����s�Y�F^,�pL��7fy��b\!��3	l�'9١����[��{y(Tt�j= f����_������5�z��
e{��R��0O��tpi���4��<ϲc����n#��ud���ou���H�tG ��{E^!!�w�`	]��'l��]�!��GIS8�Z���
��9����O��^vy��`!��L����p����-�.�Kkh[��t�a���C�$�X��l��%�;�?�^���"�;�7U�M9�BL�-�MU�e$0��U���"u�A�k�.Q��}��|B������ם"�/Ba�X)%Ŗ ����8P��'xK[��[L�P�mf�'l��6^h�m��,U��-�JO�I���ᴣ�-Q��,;hؿsrO�S��Fm:�m�p��"K�ס"��{���u�R4&����T�F\/���r�s�h�〦�����CUM�#�ajU70�N�I5�R�>qŜ�V�`��+�4>�Y�
avQ	�c��)�@#�~��b��2<��|{67fB�]�+���ӑ��=���r�N�ђ�Tdk��I���7�a	ԫ7=9�6����ͬSf:9�,��Z�E�<�1��D�e��(�9�C����㸰����(7`|p_>�G�Q�� p�Q������=i�ry*��[���l����T��C����f���h�}7,���<|٦P�BRfw����ַ���8#�󏬦�⛰�����WQ	�B]��w$׊���B���w�6���X@����ZFa|��AJ��|[RA^�[�
�0�`sr!R�"��h:�:r�0�Pti灾C�}��[�j�fbh~r!��ZD�R-�r�|�0��0hJ��ߜ(6���4���3�=��5�	��r1�0T�W��� c|b+�h|r1ݿM�+D��@/� �1�$�>�D'���l ��J‑&q�aW��Ɛ�5�綘��~�<�Z/P��ۍ=��?����D!��t��	űE�b%�*�CwĻH��k�rFU��w�=v��pm	wEc����ֿ�����)%L���]R���������c��s�1�[�|���0��g��מ���q�����O�K���%�_;�& M�;�~o�]ٱ�P�L�{;@������,���Jz��3F���[��i��Rz��~;v6��0Œ�X�OOYp!��	�D Dr�~��������x�)dd��m�n��+�� �1�K�TJ�hg�I�$���t���F֮K�*��$WJ:Q�Ղ�~�r��]�f������~m:T%@��_�*Y��`��/(��xb�+�X�����Y�G��i�KZ�L�n\�:9��{���J�瀨s��`J�I���h�; ~�x��q��]47F*-h��f�e��q�.
�!��H4�E��S��PnO�$�<�`l�4 A<�%�m~��S���`�K�������6��0U�h�Ǵq� U�դ<!Yq���$���@��F�'f���fE�@]�/�l*x$�K��Q0����������~=�"�V1������i��j��P�F�~�C�~N(y��4Q)�v�ڒ���FF�~��JX;�1a�C����q��԰�w�K�y&
�
'}���'�ű���ˢ�֏�&����חq/8��}���<�DO"�����m�
�r��0ӓ^G�)���YU!]Z������"#M���ׄM�CC,?V[[}�y-+�QTu�q;v���G�L-�ͤ��M�7b�����l��bW��;r��3Z���2��a]��\�W��P_Dt��^�������\7�~y{L��Ď3ߐ0�W�@(���hg��E&;�����F��nv_?�!�4����8|�_��!�\�����pv?j(vDx�H?�T�lS��%�%6c������Z��:6�3�f��O�H t@a������(���%e�"3�zh[�s�J���w��[��8k��=L�'��EA�. fqڣ���'(�ж��G�4�M����c��Չl pӦ_C�A����?W���ӑq�9��߬��������$3�b��v�,}�#�N$G��Z�_t��m�|����K�Ǭ����-
5_=�u��P�5F�x���� ���{��ڃ��N߶ᝐ��E��γ[$�t�:�z�2�=�4��/���~�����l���c�ק����Q�1�v��؇�պ���"^�^��Z��2�	`�'�҈�W�m��_�h�!!�8�C��(�ô�:C��-���jœ�F'�U��ů���6����Y�������uE�|$��k��S�=�!J0ݫ�ܮ(��kcB�>��S��"��� ����~�GQJG��W6~߰�*6֗���,;�\������ЎI�>�$J������
�C]��OZ�`�:���n�L~�Y���B��5FZ,*�k �`w��P�_>�����D�|I �����].�r��ܽF���lڂ�8��x�l�2=��TH^F���9|���0��4m��p8NcV��I��T��1���T���b��C*�y��M��Y"4����G*@�1��eKX'#�i&��.ɐ_Q�T�>�jZt�e=j�Q��^��M��(D�k�m���/�����9�[1/���LM�W�;�"���]�u��ݝ��.�C?��T�
�>�Mg�*���Xa�oYRu�dճR:%|J�C@�����PT���U�'��� J*>�`�E�ў.�H�h��3��:��+�`�+ i�Y�k^���]
F��Eʄ�3���z����(��|I���-�]�5�aR8���1*�}^���"oȻf�b��5��cZ#���&#��|��]��*�<�1�<A����*�}�E�g?��!�,j�V�kJ�Ku��-�Z�R�T�8\<�HۆP" � �1����eAZ":D7U�Zw ug��K��Z߃�)kH���v�M���l���R��n��9�O� qL���k�_�����M�O���CbD��ٛ�SҾKմ�9ڭ+���ڍ�j�v�c�����l��'6}cy-�+Nȡ���Ե�V�F�Mʪj)��Rt�܎��h�'*#��:�BP&K>���J�!��k��[.O'G/�l��;�4pf�V��G]F�`8�0�P����"���ޡ�>�.}��6d�A{�D*�4�ʰ�N�r�I*UՊ��(�Oi$�����[lbž.R]<��X���t���W�9R���X���o8�y��I��iD�����t�փ"Df�`L0{�j$� u���II�51n��Ng��ں�,�4Ar,�d0���ެ}�|�����'GʨI5��[�t����s�-(@���H�c�Ș�Wn�n��F��R�~Ѡi��U=Iú��I����G~NX�����
{��b��&۹Uc���P2��|%u@��1^s�Mf��<�<h���h�yG�77̐�7=�.��\��՟(Mр��=�aq��贛#��	g�p�l4�-��H��UG�r��"