��p��1#)Z`�}��ˀG�w�lC6�~�%[������1����9�mҴuc�k}r��~��]���'
o��tt���5��� jݜ�[4S�x��Yc
�⃪�ʐ�O���K|2x�9�v�ֹ��_�A� 6�h�_ǰ~�L ?	\�?_�"V�i�{��o9�^�J Ι�Z|�p��P:H+��y�u�������	��=5]9��8�4�6˥=	Y���:T߯����}r����X�u��.�-�b��[7�q�)�T��OH��d���]�G��!-q�kJ�sor�#
4��=��E��&�����뀔�r�v7� ����wG��sg����Utu�83j�Q�]^iM�2��B�#f�y��_�Y�� ��+��붹��=�Q���3<����ä��>��C�f2�3�lCL�k�qQf�@�Wy�� g�	��ZIm�X�7餯Nߖ߶�4��ů'�� ,��?��Lݞ�q�wE�_l58js��'��{��>��Z�C#�.�
?[�&�1�>W��@/9X`T���>�:�,��ٽ�=��[pZ��h��{ac�j3Ge[^�d�Zm%���Ww}����6���?ڟ��#T����D<x�����y�+�;��L3K�݅6"0�h��[�Y(5�Be��|I��͋5�a���w9���ԘiLk�U�=�����5��5��fz�����8��El���C�F�-�W�|>���.�Z�@��!�s��Dq�!�]�c6���U�by��y�c������,{�<J�\qw��$�������i�ɱ
W�$$�f緲)3�T��`���(������,��Ԛ�v�z���*G�c;߇m-_;���W�7o�����Ď��?�^��BR^�@[S��X001�V��8���ǣh�C���$21#2GJh���P��UCFV����s��F�V"��u�V�k������
�WU]�M�p499��y�b���@�"��i�أ�!!��� I��^��N~G�ʵ�{�m�u��!�=��D��s}�>�t$N?�i�����ё�Eq�F�J�8��H��Kg�y�"͸=�#���Uz��|xD�.��o��bӿ
 �� �eY+����/E2�ˮ���9��hX��y�{ez�6���]N�u��rugz�ޢ9��==���tHú_qx�=0���.���G�0=Nq���1
���8
��uH1	j�M����v�4�p$����8� F�Τ���
]��䍹���06(�9�9w	[�}&��z׼m�ToBK�*e!!��U�����-������U�k���!u�ֵ��P��M�:�{��t$�t\��H�Y8�;�L	�Q�z����6?K[[�nL�	�
қ��[|��>���;�q1Z�ҙ��0f%Ҿ����Q���;lc�韹R���q�h��
/�	�C�(�s�E�[>�2���=�ݝ�[w�����~���}�ͭB�}s��O`�[۷�s�+#����k��\r���=Mڊ�+?B�g��yB��.:B��c��	���]�w8�R��jx��z;�R����v�lx9���B�w'�Uj�|�'<_�Xa=x��{���X][��j�%�n|�KN�{@*�`Wvp�L�jlּ���V�.WP]f��a��{�){N$.DKO&����Q0j>T���g2������	C����x��)?M����L���;�"��|p�Ûٳ�7�_�^�y���<gXz��J�<��?w4��L�-�կf�ߛ&��H�/�a9*���I��������� ������/GK���5ן�1�\M�t[w&hgM��a������L�5�&�O�e��~vR3ncKlz>�ON�._DO��)�>�3�x��W���ĹD��~\r���v�w
\�`s�п�:�M��_Ms��w!?�	�������G<5�����k�3�;w��F*	f#K��`"����3mi�5h��b#V`�U"6��u8��u`��g�)*�l���eKt�z2]��z�����4���}��5���T�%���3?��Aнp
-00JL�W��}��q�F&&&�ο>_��i�-����E"�J��s�ԄS#/�%%_������E8kFby�qz�u���uD�L>�k��~��}���@�>F�X/T��� f��G�'�9�B�z=a�ur���E������b^w�6�sG�epO�A�vQfe��;���C��B�T'��#�-��`��F�7s�ey����cl{Z�d�VYuw�y�~/?S�!�
o)��1s�����t$��R�J~� ����h'p���ֶ�&V���FSX֊Y�m�D9�&9G�ϟ� ��~F�W����26�7�R���~_�/V�߶�m��$��a�����՘fU��j�����7����-��K��N.U|O%��R�}����+=_L�����E�9�x�]c�W	T�y�����"x�e�e�s����=��h9n����r�Yg'�rԵ�''_�Έf�ن�.����Ʌ��J�����7#$=.K~6��=,Y��b����ti��c����̦G���>�e?+�n�"q����+^�����੔�f��U�� S��R�׹�����O���N6��$�go\]��g�����jO����y�w�����G~�|����Ӣ9]k!L3F��Ä������h��h�X��9g׹Ʋ��w5ᴡ]�I)U3�!��sJ�Ƒ,�vB�fqX|��S#G7)��nDm��C��T&��~榝DX�t��[<6�CQD3+%\L��B3{��4�Tt��A�#��f5�*�� b��=��n��_I�%A�Q�����I���
�yb��l���B����#~�� 3F��J>]���"L�z挢�����K����C^�cE߂��Ձ;��z�v'�崴Kn��s�M�h������G;��Hl�}�uƝ��G��e�����dy�v6�+~;eQ��������e?H��r���l�z	3��l< /D���n�zZ'}�>�*�Z��x��*��H|�zߞj��־v�=[zz/B?�k1M�k�w_�zv502�޿y_?5�yN��^��?��y�}1ܽ[�H����\���1�|B��T��Z3��YC՝���ڭv�x탖�)Rww�b�cԐSo��.�y5y�F7'mߩ<^�=m��C��{�a��($q"\ӧ�׉�~��}�������55�\��0�>���:f*^vd�ڳX6�R.1|w�dA��)[]�!$4�~'���[
�[��pf_��98{�Q�G�q'!o�h��72[�?u�an[I��P�l68,(����__�x7�Jb3�O�m���ﭟA���o���XJML$�����_rJ��}�Mw(n�����-1��!�ng���*I|Z�]q��ȉu�^�6�1g�t��Ϫd_���ߚ���^��-#�

����Gƻ/S����w�!����5f+9�Ĉ����V�#�b�X���a��Bf��¡�Q��Ы�MՐP��*��H(9��:б��n6�m����C��x5<q��c��Rɂ[�$$�28q��qm��H�E���n'K��#eJƖ��U"?7_�\$�u%*o^��{�/�S�r*�-�9ˮ<4��U�S��h�9�0w��5�n��>�4w�Hwؕ����ϧ����G�ۥ�;t��?�w���1�m��~1]�0�Rԗ}�]�}�_�'��]�e�y�  l�#�U���>��?W/��mn�1�<F���NĮ�ܜ�R�r�,v80Z����FZ���d3�lnj� ���}�&^介M����>�W&�K�od��m-@5� �w=���Q���$������jK��=�j��� �j'�D�KN-	�c��\��J�r��?��}L�n.������ue݋�,�YԳ�bAV7�*��Eqј���1����MR͞l&�mk�C��ۣ;�c�1��9�*S��R�ο�٠�qM��y��wȾ��IdX��å5R�M������[��urn��|�����x����l!�0'�C�;��.Z��?P�1���k�a��T���I9,t{�c�#���)|��ohp�G��w���3{��