�x� �����. ��3�> :���z��1�w�uFH	� x0(	�p�ƙ�_gi���6�!��Ʃ����T�C&���P,*���8Jǁ0^���nw�	�����'��hX�T*�6��r��!�U��r!hH	���N/`� y&'i������/�5)��~c�p}�����!�>,�h@�@h g��D�G��z��i���%�{�GI�|@#Wt�@$@���/�;��.l<�'��=
�p:sV�`h P�0*{�R�� ��@xg!�U�Ǚli�G	��Gy�{�g�?=bH"���`�L�N�&�*��0����1S��>4�r{��Qta���l�g�x AXJ�g)�q����0f��HJc���y��2�`��p�A.n`0"1�d�Y�r�a��`|��t�A n�;����'��kqH\�aH.���t)I�z`b��g����BA�jm&԰!B�g�f&Q���H��6e�� /�c��i��A�c�#$`O�� ��21�w�BO@�}B� 
X�)�GF���
rVa�&�D0 �rNY�=&�b��P��D�x��Ȉй�b�B#\WT
郆	*� rP�P��,�`c �"�0f  x %�(w� <F���pcA�6� �"@iA�7Y�y�E�  B ,����A�	���RLK�p�H��� � �� pD��4�8���ֲ>�@ �4q�1�18��� �2� �㠞��4  �� 
A@ Q~�� � �0������/��%e���h���b�,�(�hz��91��"A(`�@� �ȣ�=�(�'(�
����(0�����t�>���2�l�_��D�0��3js���ƀ� �;X�c���0��e�� ��������n�;����w��>� 6��3j
�p �� 3��ݑc+��{���?��#�G1�4���C�"�`�8*�������c�W�q�2�����& 8�0@�I������/��XP@$+d��#�d�}D�Ts��?!�����p>�x
A$~���@P� ��>  ��P{���;I{:�� �Aκ�u�	�&N����/����xQ`�ı9�?��?Ф�.�dzh��CMi(�tN^d>�Y����י�Df���0�hi�&���E��]g/�I�X�IA@V-�Xb��= ���s@i��c��� ` 	A*EǡR�{��:G����v���8Ǡg���PD@XC$dA��@�S`�T��d�P��$ L���9�����:Ǹ���x�qx;���@�
���  �#W�t���x�T�` ���A�&��t��>L�� `H���9 �cxA�>GP� ��P��8A�����W����|z !�<���@%���pVUӱ���!�Ҁ���g��ϭ�!��	k;BeS·�V�A�ˣ��X
Q ���/F���Xza�>(�!��!�V
 �B � �F���,|�1���,��S`'�I�  � >p���Y
�2����@��Rfۓ�J@x'@�m��1���� D!��F���n�>�U��4� :G�Ðr����8���z쥐��@��p=(�"�Y��=�xEy�~�5CufB���	����
���@D�J
����D`��n��7	��z���(��#�y�C�w����
!b���kT>e��!��}Q!^Pn�:^O�-9��_c\�N�Ђa�����!Y�GS�����/$-A����e[��a�WD���2a��B�,}$8?�H�x:::�w� l  q��ihr�0{ @�8x�i7�t�R�{�
�: ��� p � 	 ��	Т�r��up� �  �S�'�؏�4�<� �e�a�aq�v��~xr�o�` X��� #�h{��� hA`
 ( I �o0|�h�!�����x��y�b�z��b�zn��r�YB� ������ ��` �%���P��R��2�2�|��K>���z�2=�(���>8  i���xqB�� X| %�;�y���m��N��v��� �	 8,p�/l'�y-�~�@젘����v2�qpa�ps8zC���" �!������ t+�[Hw� f��q�H{�� �<���� � G�/��.ș����%C\P����${����q�(v� ���- ���~`e�y�� ��p�X�8˨9�z�E�чJ�1�{� }�ܕ�}���~��� *z���3�r��6`�	�J�����	��/1�J|�;h�����9��J0Ko8��'�'��2�N�2K!��$2��e����	�	�0��.iI�% �] � @�
��x}'�y)whp��x�P⒘{� �p
��g����
��
��Y��g
�r�`�RYxz��ʨ�9�0ڐ*������qw�@pxH�y��eq?���.�� �	����h���$  ��b��S��l��np��0���*���| �X|s��c`Q�9ڇy�@�&�@'�@ �
 a��v*(p8{��y� �~� �� h|�z�?�Hi�}��/���=���؈ �.Л�bʋ� �{���(80J��}Xy,}��{�l�l~�h~�� ���� �!�� � �)� ��C��!�~�;�.�����j��4�m�pf�c��]� p�@# x��jC�z�hҀH�����\�pkx� $ ���8]��J(tX�@3H��� e��l�^�8�P�� ���$r��D�`��w:8_��[P�0���ht�o��d�-�)@ p��H�c���@��h �k�9� �-( `�KH^Pl������8� ��'��H�(H��R`�>
�U8��ꄑx����(�8���d���Xǲ؜E:�ZA�dS�@�R��0�J�!p��Z !j)� {�  �p28)�X�
��
 y�( xk�l��_�t� o��u��k�0�������'�h�!] x����0�� �E�(�p��ጊ ���h��|����H��	����jhd r��l�ܠpq���Y���� ��� 8 �>�
 ��R^��-��� ��e�����H� �"4�}�g���n,��W,x��� �(�� ���|�}!����[䈀�*'��h�����,�`x���A����G�� M� 8��u���Ť��	� k�xx�pt�`v�U��[4�:��H��5�'����x~�D�0 �wpa�J��u�ɇ��0��*�� ј����Cp &�y�a�P���8��-�X(�����9E�����۔���}V4�Y~��;�z�n��fy ��� '� ��z��\�yx,X H	�� � H��0�T 9��"B�܇ ��r`q��u�8z�"���()����
�¡��q���������*C6RA�����6������\�/A��k��{d�rK�/D��yV�E)$ ,"���FD�@���`~B}���㋁@����Q�}������t�~��oBxx <�(E`  q��P�tPF��w��k�
�(�`��a0��&������! ˰��3]��9�` �n��pw�Z{2�x�hi�e{�6��(+H�" u��.�q@yxZ�Y��n{^ ��0�x-N=����H��T�r��^[�n��T�����(H��n�q��j��v�pk�X p~����S$Xn�e'��uH`�hI��c*8��@��ȣ����\��h����l����\�j�v�i��^�}���z�X��h�0ӱ�� ���E`�f��9�4�����CؽR66l�0� }� q��a(Y�vH  ��� (m��z�Pu�W��� 0	 �#8o��x�"��� f�N�hs0z P7��!p Pr�8n�[� )�w�0�����*8{ `
(�d��[�"  h�p�oXq�hux��K�P�� �R Xlk�� ��e��e�P{ ��8*�iO�W�Xda�|�A�(/�J�h��*|M �/ ��q�*��ӈ�nT�F���@�3�Y�Kט���f�G .F���Ҫ/���t~e�,� h���/��䁘��,��]�`��H����� ��s��`�{���i�0qh�N��֨����A����x��,�ȇ�c� %�	�0п�/��R���H�u��d�`i�_� yhv��vܠm�8�u���P � ���<� @
 h�
0
&M�M!�y�vR�R�q��L�w�y-�e��y��b��f���/Z�z��0�p��#�	��:,�؇�D�Vw����E�Z�/F��?�u���)�a	D�򣉠|��	�� z�u�Hwxzr��,��T�<�x�k��{�0^�j��	�#.�x��۬" {  Lx�gHI�o�ei���8+��zI�?k��zQ���4hh*� ��0�H1�G���t�z�bw�	�(�D���,�h�s�(o���!� ���fHb�@
[W����r; pH
	���X`@������_����� ~9߯W���>RG� ��G�� ����
 �������� �  �����8 �T)S����� �S` �6�H*vy�*�gZ毧�N��ۭT�ޟN�@ Y���J�ͣ4<[��>�c0�I���m�٤��� ����+� X����|��O�Ce��l�N����G�� Hb����+���y����;M�4�H�Q+}����Ea�<T?/� �� _��0����
�?)�)�y�W�]恬u���.��`����d��)�<ͪP��� �Ʃ�V�湘h��t;����"P4 �y�g$9px�&i�}���F�����!�8 y�y�&��u��d��@|����h p x�	�� S��}�K�*��)Qf�$g��=/I����[��'����� ��0 �-�|�g��)�|�I���G�|| "��`hu*�H���;T�O�4��(��Φ?�����ɒ�)�": @J�t��1�b�Ѽe���f��d'��n����@�8�G�~�E�����x�NT�	faB���"�<G�nU�F��!�J�hZ � x/J�Fg��s�qnr�� v$��C�q�f��m�K��#��"�!0l ��$o����PA�]���l  )nC&9�q9���ʩ��8��ֻ��*��Q
�0��Ψ*L+0>���pJ�v�@�0�&�+������3s�ļ�̛�����,|��������jz��sku����r��֐�� �
�pX�!;��� t���o�1�l��{ '!��!�ѯ)t�!80��y�H ��~�����N��$`	N �0  �$S�H�(a�R�C� �qK��?���CLna�>�� �{�8���� ?�I� ���J@9�"���& h�����(����u��5�PC�����8��;Ch�9��59� 0
� 	 �
��h@H.Pw� =��&�I@6rΨ�s�ȝ�c��O,�)@��8N�8�&��	�R�Z]q8$��~(��I�'#�v���>�\(�(P7@�'` xA�,��Cw��?@� a�.��*�/#�w� �h�"T`QZ1�h���P� �K�H��^K��R* ���6G�B�w����`
 �?6v����Q h ��b�  ��~�2�b�RZ@~ d5G�cP���@�@ M���>��r@���89��2f�|��mI���\����`d��(��|�Fz��Ǡ���u���%�} �=�H�Z\�&E��d���ʖ3�bF b���!�e%�2��Jt���<��"�O�Z�-�����DO ������>�	?�&Nû�f�u&��i��� |�X.G�=D��y���lF�C��Qަ�PQ�}����H��#��`T�qi��RQ�$Ő�C|z�06 =��x�@^�X[���A�=T�.�Zǧ�P��91eA�_��i����v���;E(�c�p� `
��f ���.�ٞTJ���\	��c�c���+Ÿ��\v���p�0B�8���_�Ѿ8G��$'��P��h �����do�T,����p�B�� ��$يٴ �':����v �y>��'QZ������Y�˲��  ҤF� ��|�Gx���c��9GX �@w�a�N 9f \��$�@�
�,�P(�h��r��ϭrY�֊�cEk!��z�g�0��C$aAf3��� �0j@aR#l�q�����q�?�@�����	�� �Y�X.G�`d7��~@����mAz7@�	 �Ɛd�(�~Ǡ� @B�Z��3�� �"A�3���#��HT�(#�D�:;�x�#\sP�����kF�?��:@�`	��/�����{ ��Ol�R��(�k%��T&�̢���'
v�-N���K��ֱ8o�F��n�L-&�"G��)Ď��$M]��N�[8�b�_eDu�Ѻ��<fr)��FX ��#�$F���$C�1�
��=`���Tk���:���c�sĴ ����yyy�k����;&�X, � #�	�̈́��)� �hz #b�*$sd��b�l��3�X��Xj�P �L)�z��&@h _@@\ R @��,�`
�g����>��� K��)*�6����a������L��OK6E��0 h� ^ z�*�BM���t�@ H��¦�EÉa�B��b��e,�i�g\-H0S▂fЖ  �������١�h�|�@X�6���T��a���FF � �)������8��!����6  ��	�| fl�Ө�1P�)� R��6�^���^��`6`�`D�@ �B��j��a�P�(r�"1�ē��"r!��jA��� l��'�*!��� � \ ���H�?d�})t��|�	
 ��.�(`P  �, ���&�R��A� a�$A޳iBN�ү�Z�nH� �(P�"�Z�gB�28(V��3������.��x����<3�l�CQº,������)�-&�N�>-�e5E t`�
�H����ed����� ��ТJ�I�t#4,k8/,�e�6V�!#�����x�V�����N@T@0A����*�l�`%A� X�!�*A�P �p*�+1�B4��L�!��a�ᢦ�X�� ��c`�!�'�p�nP"�@B�&��8��A��na�!�K��@�`" �������& ��D	 � 2@�5��2A���!��Ha��� 0`r@�L�x`�L`�p� �#%	���gLh�'E�'��#�*.� u$�6.OYA!��A���A���E���\A����(�K�� �6@`P`\ 2�J�>�%����v��-��,��2�-�.I�&B�rI5Eh&E4 �&a��V�n����	���/���Zs�~@l~ ������z	`J@V��!�aF�����\ &���\1��� h� f&T��!���ak3� ��|�A���A���J"� �R�R���`*1;Nm�Of @. ��r���1�.�n�@o)'B�Q�\u��#�&(���)Y�.N�-c�/��4$�R��N�^�Rl���p&����'b��R(�1Sx0nʐb�͢|t�P�*�}&�.�-|�d�Z�Rns 8B��@
�� ��N�p�0���ҡ��|������nh !��a��a�&' �
��"  fb�*@$ J` d� @�U0�. �Td�<-B����J�������A�a���Q0�` ���!�Gb�   V�ŀ@.@��  �&f&D���$(�D*�
�,5I,+2
���/!������$���!�9�@	�`��f�p�$�&`��4.���|/"c����v��� }j�wRB}b~h��r�ڧt�B!�A�A6��!�`N��� � !sx>�j�!�xA���E��0q�za\laދa�V� �F
��`^�� /��d�Xuq�&�����������n`�@^�XM��~��,�P�G-L4��$.)�1�!�A|����*�����n���	���t�d��� �2���
v��-#�� g4�6��L(�U@)�qB�Q&��� G�a�pBdV�4.*�8�%(�e�(�4�('*�F烰�+b�gr>�Ƒ��1
�l�
�bdwB�@,�+�*1c`&��v�l�D��B��J�x @�26���X��A���a�kAġA�y���-+6ǈ��r()���d�!�� �ܤ�  r���!� ��&
 r�����c�3���`��7b�c77�&�8A���4�ta���   �	�N
��n��u���C�r&�5�c )R����������A���>�x L��j 6�n�>�T� �V���I!�!�M�v��4p��@:lOD J X`�&*M\�K������b�t�丷�VA�`qM4a�a��a�o��PJ�|��&�9� @
ۀ�<`ZU� ,ۀ@�xӤ�p�&���ɶL�I9ab�Y�I��"0��c� ���~�j�� ����B ��!�� �@LM�4Bz�E��HŠ�	 A���!2�`	 �`�a�a�!NU��`j�`�A��x ��̝��B��@��A��l F�"��a�m)dH,�� C��B��A�U��@����xF! t�p D���+�Y3ГV�"����s�(Ϲ�Q�Zcu��r�TvCqdF�,����E χ?�"h�9"�/)
Î��|�3��3e.�­(��t���b�p�<�
��/�KV 2br)�>#%-���   �
@��� b �J���� 廁���!�!�!���a���9F�-7@Q�� `L �  . @�� <e8���$c*QB* �2 ,&�������� ���!���;�F����"��`��@H �n�����$ *y#�,�+@>�#��9B>�� !��A���a������!��	
�J �]�m�@n�(x�w~#"����,� ��4-(�{0 (����j��ʯ�v0Ղ-����a������!���/|@B@�	 &��4�3}8A�A�!j��A���
@L�\ A�!�Tf��[`� (@T�.� ��02zO��F�R��D���ah���"  � �	G�D�}��cBu3��O1E�������N!�A�>��~�t����t���@b
���, 9Cꬎ(�S��!��F �  �("`8.�Q�R�qCB�������8D��k-'�C�?	*ڬc�X� ? `  ?�g� �D���8
 ~��X�J#B$p�3�?���Pw�x~?_��%� ����U�7�B�3���mM �0P�@ @-�~>/G����p�������  ����'�Y\JF~ޯO��
������Iz�T�.w+�8��������AB`� x�_�0 ��_O��"�����7 6FA��k�؍\�̗����
e����<N�ۉ��T��  $*{� (/�����z>�nW�e��q���@��" �$ @� �*�$���|���|'I�z�)�a��t����G�� 4AH��:@� ��H0 '�Q�} ��}����w�G��yg!�{�Gq�u����!�Y�n���y�˲: jp ����`h@a0J	�,��`2�iZ^;�h��`�� ���RF�<hK�����֍�ɸ
$g�D�F!ZW�����P!� Q�vg	�|���L�`�T��1�dgP)7	"�B��E�np����8�;�`8z�ŉ�h�@����xv��kO�  ���p�I�W���V
�!p(x��9�g��� �Ti�Q �.��Rt�'��v���L�@8rFQx\��XTb bzg1R?�g���  @
�!�Dv��(����y�Ƽ(HbP��hz$�����+(zZ��q�b�k	r{��2*�$8��h��%:J$~i�=#��h�����j���
�!�
�%�r%'�J|�l�\�q�zՀ�  ��8a@�5 � {���o ��pf��c�9���i�qre����潂(�f���$����d�!�h� �$� �*;���  $� PC�-zb��4R?Ӏ�k��h���q���r�;H݀ i7�T �V�( �\�@� �D�W��S�A�|��b>�iri�<~��hO��'��яA�6��h|�Q�������� �� xH�X!{�t��i&$�|�Ć ڟ �����*H�@��� c���C�aa�4��ð|A�?G������tB`9`T�b��1J�Xt��3����0w��=��S@����A��	PXQ!PGm5AZ��p���9H���u���;�Z�
�@�@pz�� BH��L����$�+W"Gh��A�2���{?2���@z7`�@v ��笗�e 
~F�A�ېY(0x�Q�y�!� �ppF x
4��b�?���c�k/!� �A�!����KHRf3��4C)�-�M�G�Lbm�C�DZ�&)���y���;M&�>Y�
\O�N;�(��XJJ������vP@ ��|��6����X�0���H$ ��&�^��m�}���M��N�z��T%F ��Tx�q�@����Q�=l � �pe`Gh�5����2(M�r�'��Q�M�<� C�b�� Ũ�Ct}���>@A!d*��P	 �r��P�Ϙ�ZA'\� !�k˔�6U�����l�*�P���p
D`�1Rʗ(s\�(�C�jq�1FX���v��>�p �d���@ ��<�@�)�� �+�:RP�����<����!���y��@R������h�$� 
�0 |
 &�im ռSNMY�' ��jQ�H�U�Ҕ�0w�Y3�M @yI�c�i�|-������� ��n�G�;����">�H��p�0��C�����3P��tp0x9����v5����X ��r��<� ���H���'Tu���2�(�7`�8��Cn�G���;��c�B
���\k��@���a�6���������7�^�A�9��7�����]�U>g�,�bK�\#��5��f+��"Dr��6MZY*n�B B|?%�"�0�4ҊGI��"��T\wZ4�!��(��E��Q���*��V>�� � ���\����e,��{�C(&	!� �f��{�Θm�!�4�X��${q�9G��#�|�`�G�&H n�: � `ӄ	D	x�4 EjCHh�oy�G� �L����F�>ް���k���1G@����Ѭ9G��?��q�Y�)`��qI#��	 (�Pc� ��ӏ4�&�"���k	9�&g������ǰ�C�A�=���C@m�A�9���ƨ�
�@ � PR�X) 8� ��
�`5 `
�9E"��*"�(.���`v��p>�l�0x��0��r��o�(|�xx��z{����� ���  �R�P����Xw��+�Pp�P|��m��q�X�   ��8 P ��@������A��؁�� ���  0^XW��t��~���?�8��k����@y�{���@�y�	��� ~�opY�y� t��x� �e�rD����0�bȪ�oX�8���� ��X�!:j�@��� �r$X����(	���(�E1��l y� ������'ȇ9z��3,h~� �گ(�K �ѰFb.&���"��m���
, ji����"��	 ����Q�`��� �8�D@ˇ�¯�q����r������2�Ȍ���(��ѵ��˹:x  v@t��Z�Y�~0r��	���[��s�
A1�(�r# �����(�	��	��	� ��w@`�XD�xq��,,��x#�8	��|�Ȧ��rɧ	��Ӎ���h�Z,�)Cؽ8I����ۄ����y+�ŇXv�@q�pi�v��k`sLJ.���yI���9AJ�P���0�
�|��ü �Y q� �����6�h�� �= i @� 8�J[w�)�����4E`�����$?���3��1aΘ������s�iHg��g��_���`� �P�� m�x��$x	�*S d�Pr�@{� ���	0kHN�0r�q 0�X`,�w��q��P�w�x�� I�X�����	0�x|Xs��\��l�(k�#�H�h~�@j��nX�+j�"��� ����f��h����	�oe�b����Xo�m�D�@z�0��@���C��A��2�kRC,���Q�KÀ�YH�	��8���L)��12��8����%���0�R-��G�&a���F��B����3�<Y������x��H��������	�

Ț�!���X	�́�,���:
Y҇�kXk��b���dE�`q��qh�H����E�(���x�p �����l �+�ܸH�8��Yπ�����@��:ל�O��gPi�c�`w�(sְ��t��4�y���  � A@�3<�h0@��5�h|����b&[ũu��:X�����a��� ��  w� u��l�{
��`}(w�y��.Y@���x����x  x ��� X ���Ȇ���`{�py u��s�q�vhy�Z#�ƃ$��� �HX�h	�3�@�����<
e��~�Q�i,<�!��` ��k���-��|!J�"������`�py�[�o���85���H" � �9�Z<�E���������^� ��w`hL]�<Ѥ  `hxrű�� )(:��O��������8��E�h���+������p	��x	 �"̇Ap�s�z�+x��B0��b�N���9��#���U��)B�c��������
�����@��S�N���,�h��虧��0�6���!��w�8o�p��~�P	�,w<�}���/x��O�=@�3�� �-k?�x_pqY�p���� ��0
/�|�hx���H&�� �j�(w�������EIan��΄���u`]pK��z�0X��.���� 0ԉ�~�z�� `���c�BM9�	��80�3�U��β��p�pכ��&[~��|�5��v��p(y��o~?�E�z;��yi*b�P��������S0,��`���X vx ������h	���]� VU��2qܚ8��[ �	�F�"iSĵ�X~��k��b��H��!��� �e��[�0Y�wh����X�u�M D��(���x�pk��{�@g`��� ����S�Hn��_��"�(5�p�Hz�Sxh�s���������  ���-�󀉶�\� h��b � ����@s�j�8Ψ�2�} ��h:��s������Xk�co� ��& ��n��\`�� `�^����
H񉴉	�i�?���rdy9؉Y�
8�ݡ�&�	�1�8��	�2��{ۚ�7���}���UFe�6�	8�ƃ�]��T�牛�q��t=�	Ǹ�9�-N��>� p��<��
���0#"u��l  r��l��f8z��s�h�xۨ H��y��=� � �(�/0�p��h � �?�����	 �  �`
�ǔ�����&p���q���i�e�`z���� �t婈a�#���@4���
��� H�p���#n3��AН�!�"
�q2�z��|0y�XsP}8w�D��p� s�[0��нӚG��ՋP�Y/)C䰋��K|b�B��ՀMh
����"8�@�9<���?�)ny�C���Wa���aK��))��Ɗl=�`�
J�E':�0�Z���Ǆ�Y�P]�Hw�&� �2�i爈u���B���[/��n㑼��`U�pwPk�=� *܇�n�(|xQqqpB�pCE�_)��� I��X�����2^d/&3ڰy w��� p�P�����h"�s��\0u�d^A)���s���/P��������ISџ��Y�y>Y����a�D=�yڣ�����%�Ӌ���P;��àꇨxL@vy 
�u:yZ�� �͗��p��92�|������    z�t�X\�O�(~
�x�(��! s@�gX�z � H4��xr�� yZ�țȁz|@�����@ R��g��w8Z�tH����$� ��&�8(9����;�����ᚈiHB�*��Y���(������ԫ�
�i�2˞����</S��n���:�Og{���u��o����z��ow����}�_� �`�( ���0� ��P0��D� ����� � @P G�S�@ $p � 
���� #��U?�*%*=i�(@7�U�9��b-Ά��6��`TM��q>����J������yC �Q<A)-�B���g�8P@�d�,%�l6}��@��p　�� @ �c���h,؂K>�.�#E��t��������Ĭ$�h:�� ��x G��b���p a�� `�"b&Y|P�G�� "�������h �j*����y��������Z;��� ���������v�Qʌ��0}�����j|�+�)�2��Z�~����� �|N���J������r�V����4 j:��E�����0쪺���sA 3��?��,��G*����1��X�2��P����B� �u�a�~��f&�{�Y�kg�sI��G�����&�!�@����"�!���‽��s(� 0 	  *Zq� �Ƨ����w@�g�I�i������i���{N�2 ���8n�� ��
 x,��!�."��/��t��G�,~�
��'�P~����Ȳi��(��~e��~��q�q��u�H^�v�gi�~����y��ܘ}H,���G���+�<��P^�H	�.���,��n�� $��Ч��"�'(�(0���Əc�9��X+(��6�K�j��P�Դ�U�Er�������R�YV_Ǟ~��P�8�@T {�|)Α�|��C��Dg�(@sgQNe��!�xQ'�2
�ڐ g�ǡ�r���4�B�V6�� v���z�nZ読H���yt��JqOEH��!�8G0� $��>	��@����iBc�|A�=�������?�K,����B��P�6q���t�א�8E�!<'�e
�cNk�}�Qiu�q#$R�?K�Q@R�P ���l���=���c�q 1�9 �J��v<=ܘE`Ba��
�nd�=��.?���H!n0G8���i��>��L����::�p�C�r?�hR��� :�:��$�v>���ce�;��PJi4#|q�<��!C�|��4B�X���. JQK�^�@��	IFh�Өw@�
+"D��}�<SٸE�E��2��Y(�H���f6��`2�l����Ǣ�(�0}�a�=���@|��~���IW�4 Uv@0	b���@�J�M#��&����!X'�����\��(���8tV��5D���y>\.-E
� X�F��"�Z�A�3��`�� \#��C�}���[�(�Xr�2�h�x�(`8����M
7� �xn����88�B�j��=B`=��#�@ T#�{'c���Q
��7G(+ �c Q�3 ���{�����rc��� �C� �1�<��I�T��0������N��6b�i��$3��C ����J2-LS�<�4F�Q�?$(�(S���P�"'��6��Q�FOt@��%
Q�"A 6��B��<q��k�N�S��H��f�
�?Q��!f���0J�9��(�Ǚ�~)#�(�J�r�{��K�*�T-�Z
�  an�Wz7@ ��͢Q�:G �#tw�8G��9�m���1�`��� ?���@Hp2S�n-Mi�� �  ���:�є;��� �? ��qA�>P����[v`�/�j  �	  h
�@4�� � �Yi}��(�\�.m�ނ4��: ,�@����޾d0�k� ��1��|��<G���tP1�;����{��?�h��t���ؑ!ӂ����@� �� P0�8` ���)���ȳSg*QѶK���e��G\�.)䨹yH��\���D��ӹ�%����0X�b������` �<�F �a�� 5����!�)�@(-�FGp��d��v3�x��o 8@P�C�d!�EG�B \D`k�Ԋ�2��Q��j0I��' ���)��� T9=�t��@r���,Ə��?Gp�l�����?2�� �3������g)=�#4��J+)����ƍ�S`�m�@�����v.7��Gv��jKCL4 �:S@jL�Gg��G��`'��Ue礩3��ވ��]L�������]��u��r<x���z 0 `\
����,a�����h��X` �`�@���MJVeg��F���� @PH2G!����������t �
 N�  �@��6�h��ns�<Q�:���)�f�)��p� �\I��\N+�c�e�^O�v�(٭��(D$bW��Wư#ρM~eb�d�H�,���FxGD<#�<I��)d�~�һ�L��@ �V�>.����G(��I�>p!�.�&LJD���IȒ$�#a���!�!f��`, �` �<���-�{` O
 
A|b  ��`@��! ��
`��� R��V�����z@`~ �h��.\�y�@C��aja��� 4@\�6�a����*t��)���. �D�@�!�`.o J F!��v��`@r	�x��!d�����"��b�G��)�)d<(�D�I������:���O��$�CH�G�C���E&D O�J�VW︄�BG  @� E��=h�"�&Т,�j+�|*��P�C�BĀKel�Mh�Fh��DM��W�BCĬFE�l`�  ��j(��`��H`\@ beDT���zA�!��A���!�\�JZ'����4 `R b��> n�*�&HE��~  w�(� ���P~�e�
p-!���!��� ���%�Wӈ, C@D��b b�&�^#�. .'B�#e�/I!+�H�P�"s(�ee(�c���B➭���|�d�Enx"��\��Ki`k�"�������F�����//����j(�@ f� "x+��r
+��,�d�ⴣ� F/o'��>K�4*OL��|����Ƞ#��khP�0���#O��b�����Az�na� x�. ��\P�!�\�4Ŵ D� �e��O2r�+�>��A��a��>7�V �vo"���>`�`\��ZH8}��(�L�C��f\��#'�No���(W���8a�a�� &@@��>:A�	���Q!��Z��Z��� �4o��\)Lp�����Ό�M��F���:D�S-��l�<\�D��O�*� D)$��v����(�`x
J�U�FfZG븄� ��'�I��W)��� a�|�$A����4�� @	���8�A�ar����`   ���:�$H"� �`Cb�#���Ԅn"����r�f!�!��D�`��l-� ���s�ԉc,F�"�G�,E�  $�>�a��´Ԡ
��O�CjC;�6cfx�dr�ĸۡ�j�W������s�����ND��R�
NH�)Vm�@��)l���]B� �:�r���"�"�l�4-_v��/h^�'�Mic&,4����� a���a�!����� ���-���A��� @J��8A|��!��d 6�|m AL��� p�R��$�aXA�EX���@�p �"琠��9���A�@�*�`fa��A���$`���#�l�  d� �I� �f	�x Ϝ�r�L @8 l z���L�A�"H[G*I�����o�d)7~��M(R(��DGF�4.�bP�X'�>(̀�b����d��% s0�D��ٌ��W�\J�,GjF­v����gI�)� F��I�-�~C�\�LQyĀDDxB��\��\�|.�~�  �dL`6��`R��`s�D[ED��!��!���9�����sa�VD~ !�٦�  X��. `*�`X�@g �
��OB�[@(S�$�%�rp~��(  �H������!��.�!�����F�ZW� �: ��`fJ�l�,AĲ���a�k�Fs�+����r)�F(��D#�H�#%�GK�g���J~�6�����c���՜.�
�)Υ��+D�f��
��2��ܫx,*+Q",��N�)��8��ea�G��g�`Qb�'�$��Q(��GLb�\�`\�8kdV*��J���� !p ��`��\�$�/r��D��8Mwp� ����An�޵��-BkoF/�ax�$``d��f@@E��І G��`"�\b�N�bx�8H��Z��Oͼ1<Tf&�Tp�|�(� ��L�a�(��)B�I$Pt<I˸�C�.����eC�I�ơ��N�gv�$�Җ�i,�^��  �"<D5���a� �* !�2a���9��[D�+"�I� y�I����J�4���v�� ��jA!�a�@D@
���p�6m ��!hA���"J ��@L��g�ʷ�:`�g��,+���E"���J�4����������� �	�V� ѢO-g>rx�vD��i�F��#�Iob8� h�� 
�����H.:��$��m�e6⾆���`�db���-&L��ؠ�c:I ��VA붣��B���l��\���fDȥ�:)�v-Q&���E'.*�*�bN�\*g3u���:��I��.Dģ �n��!t!q�$� @t B!����f`J�@8�!��� M� �@:[A�r!<��z@�� 4`AP�lA�p> ~ :�l�2�t [o#�$��ŅA\���\ *�$ a���0�?H��Z  6�
`^�w���fv�8 ����v@`L`���� �������b^�E-�Ŏ)��fI�M��0�FDU��n0�g;JG=�iq�ݐ��-�V�  "{��5ɽ�l*F+�C�C��5�."�B��,pK��s�T=� =���G��Ă�0D����Ef�6�0@��T	�d  ZC�A��A�������C���)S5@'9�Oa�` ,  �J� A�� �� �P�� >�  � �}� �� PD 	  P$R,  ��|q��F^�@i��h���绥� p;�g+�����Q��Jl5C@P|2���� `@4�A���U�� �/���.~�_�������߀�W��d� �_��L��k�̟��u�^�|��Z:�}�n80����Tn8��-�a�����P@D��P0$݀� �h�j�W����+�þo�s���}�_�k���~�<�G�Q�Q?�Y��3u�"�[� ���(|� ~�G��n�a�v�A�y��Є�D�A�  �z`��30�"�����Is6 9�� x�Y(_���v����X���4���T�gI�t� ��c(V9��} ��  b(}�R�� ��J^ͥ��d� 9�{�͘���x���{��*��H&���~���@�p����t��h� �/.�n�.��5�V�q:�SU�W>�KV�O�k_F�H�Z�` * �}�gz�w��Xz�`��S䶪  4�eQ7ճs13��{zհ)��������G�,^�e)�{F��  � �"|�@�рF��v�幰g�gb>��L;�a z������%�
ҳn������`'! bfY�y�'y�����,!�\W��� ��aT.+��:.	�\8�D�@N��k�8F����|/g�z��ٷ��� ϴ����sZ�5��� �`���l�~Z9�R��Ȣ��a�}�{�y�'��|Q�}����|.G��5��"U>Mκ]y����A��k���\��q�AzU���>�Nz��&�Z�Wꊈ� n3gz�gš�YG��| a�^�
xG��s`"���H0��� 3q����(0,?�P��\Tp �ph��*7E���k �>A�4 � ���yO��z�2 x���j1z4���� 6�p��pm�!�[ɉ�C�ۏ�2 H`Tv��8G(����jG��b�Y�����4	���,����q&���%����0֊��)괕��0T��$P��îES��#&�7*�\$�&l�J�*aL)/4ʵw�@c@x@0�
���zC��v�u��t�H��'B�_O��&Fb%���$�S�u'�agR_S:t/Ȝ��sl}2�-�Y�l� WAP6 &�� ���� x�@r�q�;��� #Hs���?��_��&��� #����@ pr �'���rdH�I3Q�,S#K�b��>�U�mDpx��6�h��i��9�X�#�kTQ���Y� d p	�0;�
��" x J� e��I���l�\�C���/>政�����g1��w�ƯdJg"��r���_S��-gD�� 
�0�� �X �,
�0` �$
8u� �C� ̪H�BFe4�]�Ӧ�Z��0&4{�q� �����q�?���2ñ�76��5h0�� }ф�/i��;���c�Q���6F���(�`�	��e� |�0 ;�y)%�h��\�dM��uT!.G��#���Z�hG D�9�h�B#�]���G��1 HA`b�� xv�,>	Zj� J�j���U���JSڀ"m@ ��7� �`DD pC�{�cG����p�Ҥ
�Pz�y���љE��MJjYd05�IW�H�+�R�n��<}@ ? f'�{Ǜ?����@�+� j@<K�X '0�����?��������X�dmV�V{ �BD]���4��@� ��X�D �@8�yj6E��c�z���A ��%�'��H��"����&���CDw�|<!��àw�0B�M4$P���*?��Q�p�˦\FX�D�IP9 M��'cL��#ǌv��;S��eD��=�P	�~}��ѭ%e�D��TjO1�#�  q@I� �K� �� ���-��5��@��a�=G��Jc�u�����X�ED�:�ҢXJ�S5R�����e@��# �߬�Q����\�swMd�ۧH^7F��� ]��<�4� P@���`ρ�4'Üx�₆,XK	��@5F(��r�� � n!0+�4��c<x�����	 � �VȎ$�`�fǸ�Ci�q� � ���;F���8�D?�X��`�G� �cr� J`3`z�`d��f�m�x  �jh��KX�r�ٯ��������IÉ���Yk
]�$z`�b����e&*�
_i�A����9 /���1�]�����?�`�q��ʹa����WP���YT"ZE�I`��ًqV�H��p�x�%�Ɉ�����Њ�`�Re�`�x~��7�3�#� ��	y�pu�r�q�k�ht�h� z�f����Q���� ��� �B�P (���p� ��ʎ��0�rI�  z���� H��Q��8�|��w�� i��d@i��z���w�m�Kq���X� ⧁� (����r8 :� � ���ʰ��뱚�A��	�- ,.Q^��+i�&�}����z�B
�����F��������,�
!� `�� ��p�ӛ��iw��z�ԇ�w�P���ڙ������� � ������_�y��޸�z�!L}��q��z�H�������:��ĉ�R���⁢�u�Y w�dxu`}���6�-(��˝Yʭ\��(�!�]�j�t�xZx^0�r�X`�� ���`pxh]�Pp�h|��.���+�YEH{�,YL��B�/�KM���`%�՞�y��� 8��s�t��x��
�����ÁH)8�hy��>���:h�����Q����UNZ`�ӳ�9�-So���G�������u�0���z�'huX�m[���A��w��u����r�yƹ`�ߒ����n8I��v�i��p(x���H'@0����ǀQoHu��_0rhY��r�@z� �A���E�q���&� �����s��q�X]��W�h �w��`"�)` ��h#Șؖ�|���
�Ѷ� 4� @�8 �3�����y�3*�u�v��Ӈ -���* ~�(��׎���RΌ/�f�4|�
ۯs���	P�TX~ @x C耈����� �� ��J��rA�|�#���sU�r���.%��1��ؑH ��.��X��Q�9��&C��G�;��c���GS-�  j����]0l�PH� 0%�q�;Z�
��@�X����x|��H8�h�P��d��~�p-�`1P��r� T��g��kx��	�C�� ��	����s A�M�p�@d��[�~��{�"~��w#Ps��؀	3��~�rс  ��p����!�x	�h}�^�X_Hz 8( ���`c(ZCf�x�U%��G��?�8��I�>"eA8�$��SjU$�8�\��zN�,YE�������$"g�W�͡���D�����7+�XJX�b]/�4X��$������Tk����9�H���4	z���VBX���	��� �*���@� ��Hu�����w q�xexp~�q�j0~�H{ �����t�x ��ǀ�>�H�`��wŜ�� )`
	@>�I�����Y	��w�1��ipv�l�ڡ�o�@o�*k��o  �x�8��p �ƉH�h	�p �Z)��G����.˨�k� �ҋtw�K���(�ʪNjh��V� Y�Ӫ�����X
���G�0|F
�U����Ԯ��s��z�u�\����x���獁NV�~f�x���8��in�c�	���0엀ˇ�$�p�x�~�p��{����*m�}��/��^��v�Xl�S�uYy���h
 5�n�|�z*Q�Y�u�aх�pPH�u4� ��"�	0b�(��r��^�Hw�f� x�8��.�x*a��)����81�Ar�&�ֱ�=މ�-iɹ8 h��v�`opvx��a�3�`����x�驊B�������2��+�:*�����1�f��%UՑ]g�K��	 �Ȋ� |�Pw�x f{x�9pp��o�Hܸ�D���E�����i�C)�P  ��z�J��q _��t1�P��(P�0�a�������Ua@o�z��x9����&)c"듇�ѭ# �~�hk��H�yPd��u�P{x|k�`# �"#�ޝ����㉨怈 p�[��O���pw�Pn� k @{�0�xTxx��}���N�n�D�8��i���U	x��i�ہ�u�"����ˑo��} 8πPz�f� ����&�� �6��ޚ	zFJ�td�-�IH};$���ɽ���J�Y�d���N"[��i:VQ���hu#@b�Y��p�~V�  0�M��v
CA��� 	D P p]�Py � ��y�O��n<(z�H @#�y��N�Xf t P"�@ ������f�тR]Ac(]�po�����h�@v]�X�(��( �9�@ـ�H!�Өv�j��`���' �(z�`��e�PZ���k����5�U��\!�Bb`���$�h%�z`�@Wp��&��^8��*%%�CiW�PŜo&�8���̌��r��z��H���eM(�h,qI�&��}��b�8�19k�P�J�x����@ ` 8 ����8�P?��B�� u����ۇXe8v"�|��s�� `������ra��� !h ���p�`�i�-0����n�	�@	�zʭ��&���o��܆��`l_%� t���I{	H� ��� M  =��*� h*߹���.�B
��jlVT�x�U�;ϒ�C�ʊ���p�y[��8��c(,�����$�O�;����se[,��zu���4s��߇�����ᾎ�M0��L`�p��3���u����	 �� ��t�B �[��єm?��q��y������!]����/�&W�w�pb�w�H^Xm�{��
�@���h6�`
 ��� z���   ?��0 x<�MG�=j�fFaX����@h"�w<�-V��^�v5[�Xh �D��� X y;��K� � @ :M(��_��� ���� �>�/���A�W����q����`8�� p0(�{:��8����_��i��G&���6RT�Ca�*��� ���2�S�_�jx��ڪ�l�n�|���#���
�@�g�)��}�_ 7� P�a�`v~�6� #����5[G�9� ��@ �|�t��G��mǡ�{��8$(�A(h�@�����@;^��S�晄d1+�'d0��Gq� ��� r"|橦u��Q�_gɼq�@#j@��%A�b��xB�Q��!2���� P� `6�  � H~���y��	�n�i��G:"{�'���*�| !�3x����ă���~)@#l�B��=�a��! B6(r����ة��􆪈M2跀
�z*g����@ �H� 0	�G������y�'�Px��E�v)Ǫ���s1D4T✨7L���Д~�L�b��H����� ���  ���hEy\p�����0���w��q�~�p� @�fA�w��p���|!�!�z���Q�g@4�����`�i|]���	bH4a� �,� ����� !�d��i�`�4�AX u��1�s��k*�A��H������@0N�%�fj�(�l�&!0g�E�y�g���:���H�ʇ��j"~�Wj�5�Z*[�s"ѩj��� kyA!�V�?����v�+]��!my�c�
�^��
�L��P;l��Ӫһ̇�ʄ�AQ
ߪ��4�0�O���HR��6ͪ��+
hL���\�PS�%k��>����	C�{��B�j�* �I	  x� ;�� ��j���4Ơ�#�~�q�?F��\%��s�BǠ��, �& A` `�� H@0. L�0D
9�!���dA @e3�lUJYJ��Ð�2Cc �C�h!�3ǐ���u!�50���p��DL� k��h	z%t� 2��.�|��R�U�{ŝXW+%R�I*��ǔ�J�^��3�=P�
@ ��P � | ��$fIQ�#�{���;ǰ�c�x��=�rD*@w����)�!c��N �*�+1D��dS��9y�<�q��
�8��~M��
`$�P �H� ��@ c�0��?�b�\~!�Z�c,ˤ�Jx>�x��v�!�+���cv���? � aP$�(	xw���!K!)���:�����^���8G�,�0�6
@�
�Hŕ�;�P���Y��7�8�@dL (/���r�c��Pv��(��xJp�u�TѾ���HYn^#�w��:Gxt�
�@
�
_ �(�1�;G�BI\ȮH�B��b=��1����J���9r.�D��MF������' �A�=G��k 
=Ǡ�#�9"w]��H�p�6u�Rn��)3e�@ k  Dh�!-�p�� y�P&�@Q	 �!��D��u��מ�8��h���a�R,����P.C((��	���D�p�q
q�=�P�Ðs�@d��=	a� V �FH����  2�re�� ��  ��?���İl�1�6�e�7C�).`
��Ә4�i�*+J��3�ER���fOP�,��?W\{A]�H��e�^!�Ǻ�R�	,�_���k�� +@$?�H�T 0 ^� ,C��3l<�0��el�(�zdWiN+��� s��2`��V��^C<$<t�q�1���a�A� �����( �<+"�� ���
�X��	���@�p�H��Cr��@9�H!�:8@z��°U� <��"��aFC�P��`�#dA���00�Y����5ǘ��J:.9`  "����!�>G̹� @;Fx��g�	�`I
��o��0p�g� pK��Ƅ�C2��ݼ��Ak�B���{���Ԯ�	"*�ùSƻJ��'3�����V���7F��� A�Y`���GUu=��J�Q+\�<cQHU�'/]���<!�?�;��S$��wy��<����W5^���E�i�rvq��X�P4AL4�``�,~� |C!�7� ���t1�2�8�C�nB��GJ� ����ҵsMz�@\ ��0 `��PX ���Lql�X  "� h��b�*��+a�)b� �.b�A�a��A�!� O�������wI,����* @�`�XB"��� ,�� +ð���S,4B��������\)(6���F)�    @��D @ b� ��.L������ ���������"��3���x,D�,#��<�V<k���[´�h�J�9x!'�8�h!�Թ�)A�
����4`$	� ����ɂ!�A����3��:��)��:'}��MC��������~A�A��� ��	�>���*0�"0�� (f���!�j�!�������,��Tg�!j �A\gA|� �Z�$ ���,28����^;�</���5�r#N|
��� ����h��!ң�@: $,�+�:!�2�� ��I�\��i�)i�)���IĜg�7GBub�w�j*C_(��5��lA��
��K� @Bd�� +.�Q��KB�GH+�D�EC�x���8��A�Ap�^2��� @��:	 ��L *PC(���!C8� �a���!Ja�Ī�

���d3�����JA�!�a��˘�V  j ,��N�X �k0r��3	�l� ��8��v2��P�A� ���� 
�8�C����U��Qµ'K�x�&3�vQ�l}��7I�*'����r��}�=�^���wrċ��x��*������S*-EQ
!��4���*��/��6�'�h!��2$$2��u��sB�\��ROBt����9b$*��A���ar������T F���Y%�C`H��& ������<�, �`$i!����`$
 � l������@"�� "��  j�)�)���"!�a�z*��V$h������-����0 @,� >a��� �d�H ��f�f�8 �$��^��O�|�b��o1�@G���Vǂ�Q#&�� =�t�/j�$2�ED��Uq�R,S���� w��r���&���T.�0�ޕ�,�\",l�*�lsh
7"�*��Z��v�.T�U�l1�&�%6�kN�B�2�D+#j3�.��=@|��<�=G���S2� �l	@:
 ��B�\��8E���H�����A�A�����
L㺏g� !��$� 5T   �YH�R 0n�2�G�-"�"� ���d~��U���c�*�fà A�����T�!���A��� ��
Q�DL`���F>B�$��2`�b�j�}�^���U�7Cj���~��Qâ<��
"�9���W �m��F���A� a��&�� r�<�b� �X|�8���<�;¤)'**/�K��$�vBr3�	@b��ÔCT8��3�@ a�  �.@,��G�� ]�!�A���P1w��#&M�b����fa�a�S,� @�@6`��L� �KGua�!��D�A�I ��	 ,	����P��S%� Ma�!���A�0� `f`$ �`rP��乀CA�9c:�A� a��wS�����{a/6*T*���a��� 2�I��p���P����mP!�P75�,#P]'�1�"u^���[��MB�u����\  *�+l��"1`/9c]p��l��;	<�c�r�4��tKR9"e8��M���������!���`` ��D�+��D�0�#�2��4IL���tA�!^���@H�`��`$AfA�!��R=+�< �f �	 J UH�$/�������x�'< ���!��������a���#�"bR�v��J��� Q	@�ojv�V)G�',�=C��Ht�3�)�V�CP:#.�5��BU�BwKW|  )~O�� ���������.,����B�+6��`����;TLT��R��t��J�GAxa�!��C@pW��EpA�ˤ 4 �$`
�u�$`@�D�2!�l@Ad�A���@��!����8�����|`j P�X��	q:B� x�ǀk��a`ܨ`h�� !�����zǌU�   ,``6�"a�����@_7�l��G�����@R�(� ��O�<�Ln �P��EXt2��t'*]��=K�KEE