۰p\�gu�^P�d���W��$���VF+[������`�'H�M? ��xo @,�u/d�{A�Q�e�L�zi
jݦcl֌h����ZX�q�z{�� ������t��z*|�(����!�:o�aU��7���H�"�ڲ����?���ƃ�J�Էa�Q]��ô���~�1���Q�ʁ!��9�/�ɉ��j0���������gb-��y��`��È�$��O w��!h��@,l:�cV�4a�E�f�7�OB��Nʴ�����G�<�=�I�a��b��� �qt�����»ၿ?)�b��IH	X)w@[��*��|w���X-�nv���ំ��27l�/�x������.�T��dx���ò��U�8�y�0jz���oպXZ�����۬4g6ɗ���'ٗ���W�i�x���ȴ�� *_���1q�؜G$p�Œ?5��vF�#1��f�Tثk�}&Ck�#ݮ�c2!7qT�&ĆW����!φGz�ه$�#"eZ�"�����lɅx�������Ă��,&]�����SHV[	�h��xe'T����Dcq&��إ%���/5ވ�bku��.�+6p��S�ϣ�a�'��~I?Z�W��a!�j���3��cKs<cPp!�O DE�ih�����:Vpk���;�'X��f%�:"�,%�-�8nNh����*�&��d�u�!}��늺�D���#���#|p���t>t��Km�
�YG�1��WaO{�ap���l|�S��X�Cg��z�|��������.�jq��_}�����=s4�X0�YIT��o��GHE0�L�y���@� u[��,��j��Y�|��B�!v�c�$��^1���I��5`���;:4W�/�W%��[�*��Y�8c?;� �+<�<�	XLg����Iӝ�#Īu'@�h	�Z�+�3ڌ�ϗ�K�>!��7�r�	n����t�A呒h�����Ǖ$�*'�G����GЋ��{k��
j��4iѸ��OI	6̏3*_��Z4��k��B���3s��!{	ݻqǗ�D�U�֫����%����q��G�V��c}����s&���s��U����ƞA��u��!�W`�j�2�9a��5#�s�6�Ya����IzcaE�Uhf���-AWu_ҚQ_�!���@�C�A�"]���9Tn!RΝv�t��d0 ��Ns�r�D3uvG�Eծà��l�9*���h�W�ˏ_�����7�:�ӌ���R��:?/�i?*ȃQ��K+���f�Z3�ǐ�H	�Nh��L�ذ���>�?����Bw4
@����V)b�W�Se�ܢ`�o�����n2 Hx�ơv2�b����k3��0J�ю��e�9&���r.��pI��3��`,�c��#w�~�0eʹ��Z�hc�8JUgaiW"�P���Kʎ���\|b�
~��g��(?؃�f�G\i~,ܘ��R�NX촩Փ���;���8�R�_}��T��@��r~1��H�� �=APun��|YQ�ezY���0o\>��5��Pa�L\�L���GO�\78ί����\,A���
��vw4e�D�`S����a	�G1�MGX6���~M��5��qZ�K++���]ϭ	@��r���
VwNr;O�����P1��9ʫ{�x����
���7�I�uG�m� `/�p����,�H�)�8hK�!�d�N��UT������L2|pd�C������k ���ps�4�ۊk���aC�P����/��V��~IE�-��:f�#���V䞙�Pe���tF����T���SsK<*�펑�j���V�k|�ֹ�ȸ�ս!�>�
`?���4�XAb-�_!Ω7DO�ο��lΡ/r��4 �����%t��v�V�y&�)ތ�dA'rBU����OwfSt����O�Aa'���b�AS���u���Ԯ���U*uPv5�|�Z:�v�r>��d�q��諾+��kBP�NK�47�w�j�qr<��q�=�(���հ@O�M��R�&�o|aB�ɥ�;�4���*���"�c=��rӃ���p�z����P؋��3���.��%�k���K~2p@�H3�u���ҫ����ͤ���ZDy�����Mi���QÊ�!3'�^㣗��L+�(�;���DS`}�9�ל�G������������c����C��A�ײf�`҂��D=�0�����w�#}���B�lMݣЦ�L��)���U<��!��L�Tb��3�������yg���B,��� ���g*�mG��F|8uޖ��䩻-�<w�#�����栬p|�J��nz�)/3�q�II�/�0q�}P�Va�ҵ�� :v豠�JN�S�q�;!N��������r�7������	�pI���}��M���jB)���n������+`��[�����:SX��E�f'�뛿,��G�(�4�j�֪�Mg��7´�������)�����u�!Z�=�q@���Bd����> ��c�ۋf��H�i����7�#��a+�>C�iCB�<�'��`�~��
��.�)� �	���ǔ �T�	���X\h�C����v�p����}� p~�6P�G��+|vh����M�4�Z�̏�R�v�pc0���8�2PA�/JYˢu�n����$ɭSå������zhc�@�R]������+ut��^u���c�C��HDu�O ~�#bA0|_�4�$i�;0,�ӣ�_�|-�ZS��I71���9|ǃߔ\�8�R�v�怜TU�[9�q��6f��WDP}�'47����:xqc�O�;�4�K��-��O��[�z��z�P+�P�*���҉�k�V/M4�0�x�;%2�?m%�����&��@�29���WU�T���Oa** �ø	&fE�F��4'�BS8�K*#QX��)�_�c��O�3C�{�VB�=�$����!~ڤ;l����R$L�U ��Z*Bh�I)��XqI� z��<6����z �L�V�<O��'^<��~�>��\�;X�J����d��ӧ ^��L7�m~i2Kw�d�k$��EC��O�J5�̓����C���ؤ�0��;,\b�.����Xn&0L,�q���.���|C�������o%��B{�'a�?g$��cMn{�t�zy~��-P֝o�	7Uc��G����m�(+.0���;M�v��6x�%�u;�Wb�E�d���2���\Ӳ��+8���B?���'����lw�l����g͵�!Չ1�1k�k�wD-�%<-di��hy��g	7!}��;��Lx"��E􇐤d�UV-�Jt���]�I�
�MH駎wF"Bt�5��B:
��iy>�qM0&k/\K�Ҿ�����jfz���sI�)���\���:�y~�h�^�^��ܩ"L߲�<<�S�4H��{���&�C��pAZĜ��&�����`?"0g!1�s��4�y��}V
�S"$gp��߱ò"�HnN6�Q̑N�F��P"�/㾿��f����#�5g���N�r$}l���"4J�C#�A�)Y2L��o��{B�o���Tg4J��U�}y�_��Nk�i�Ɗ��B.,�4J�u�A���lg��I��4�|�Xryt^/M���1b���D�b�mA�E�?�`�W6�1�1)��뒩�<΋e#U����D�Ѫ:{#e�X��d�;f4�_K�5�nu��o�*@�e�\֫]����4j$�� �B����"1�@�/*�����0ݵB��A���	@��I���b�B�#F������B�0׬���rK.k#E�t"jz�-�ٴ-C�w%��v��ô�-�¿���A�։F��Ɣ� �3X����B ����"'Y�!�
{�P�J3`��%��0��vog��@s�G����!�Q�@�[�3|�H�[�!�E�SJ�8N����q.�[i��?v�Bl����n0Bl��I���6oO@kI����$��M[$����
!�@n��Y�Ѿ��JӺw�Lz���I{p'~e�{��|q�,�o�KSi�Rn�A�ڕ��C�t�c��!��r6`F��Ha�PLn������=q�&_��d�O�q��A�E����M	��3�+,A�w��vrci��8y�*���_��m� ����ZMV� "l�|0�*�D��Go�R��B����ȣ��E�ܮڟ���8�N�]�ˢ���N�Fe��
K- ���U��`��%������`x�dL2��1����#�c7�Ã�����A������[fT��aT�	��v���[�6�k=�BRE\�;ur����x��ƶ@%gaU!��jM�ra}�¶o�q��̿f-���M�eN��R׶Ø?���;_���F�Ym5�ЋJ�%�2�PLMY!ň�'> �Gh���!n�t��'�ːU�E�E֧EB�B�%f���~x�ǚD�D9��x�nh�i9 HM���z��"!�\��f�K��γ�Fch���V ��߇��x$��b@�?K e("��~��O#�M���uj_�7��*�7�q�T�t�'f�~s��6������M�Ð����9񷟡$� ��d��!f׉#���L�TR��E��R�4B�f-"h��&;v����E5��}xw���<����U��,7ШdłY6���''E��I�|�SU�|�����}��釉����dI���	BkC'`u��� �e��ָ��rC������OM���Ct�ජ�����O�P���Ž��{��nv����h�b�?��C��ee�tR˓�߲㔌W��3�c%���K�`�*�W�e�WBӗ����b�/۝���Z�3:��	�M��5��%�p�B�v�C���~Gd���rI�x��R����B�q�0jh������2
J^�R�Jr�ޠ�
9#E+g��W��B�Q�*��m��f�	�~qt�����[
�R�ڋ�䉄j�9�r�ό���QM-8$��3m� �8D� +5����9��O���{�Q��WU�����*��8n����m�����q���L������7e >f��12Bܲ���t���@��:���q���	��ڔ�.�Af3�B_�TO�Pӯ�YV�}!X�AleD$R�V����c��:��6�PRP��N�d�hT��Ⱦ�ISq�#I�"�W:ׂ 5(�:n��=��3Ө�DD�UޭF�'�W��BP&�ϵ�6�w�t��DOH����4��c�<Elc�Q۫��;us�܍��wĩ�޽u����#�@�R�6������;��P�l��
���GV/�/&4J��JaF��]u`)0d�Qf���J����m�Bd 3U@���zZ���'��N����D�>��VI{�Be��7��Gk�����,A��~�s�
�>j��i������������@��dF�#2OV�j?��Ea�P�5�
�&A�<_��:
�_���/�Wlz��w�9���
�� C�lz�0/	zya��8����`�4�O٠�%�G��2*�BL��p��ف���3��2A!�����޹���=�*5Q�6��E�yX,bic�&?��X}�E�V�m���zd]����;��t���w���[2�
�0^�������DFڠ0��IaZ���̌^���ZT�O�'-��un �P��� W�;7i��.S
Փ�&7�o}�-A��l��r-�<h��Us,���-�ʪOg-��f�&)C1szSl��|Mc{;�������֫ǵ�a��%��A|j��@b�Ϋ;^IkP���`Q �z6�lJ�d{7ur.�ź�� �qi!�Ʈ�����?���4e����.;l�_0!���������\�Սy�	|텸�o���y�>4R�8�� ����z"�����Ԩ �;�5=dh�H��a��Y���(vgs+�QW�3L�*�O�JRzu5�눱��7P���̊p`3����״y7�i����V7__�(�����c͞R�E���/�Ri�ʢ����F��$�FlQ@����M��������Vj�H{_��1~7JKeHZ8J?�1ǆM��wl��NO5c2�=�3ҋB��z�#�Qп����paf(����A�?�������$�{l�Օ%۞�����7�0]^��1)���}�6"��`]�Vd�m�PdDa�+n��$����T[tr3�1�GF�,��� ^d�{�O��M�sP 8`�EE���2�Gd����$lI�#���];ٵqHJ|h��Qy#��S`X��L��H<�u|�X�,��O(N����B;�a@�Dm�6-�G�B�<�= ��S�p#Go�qw�M�d8����kU�������$����LR)c��p�����{Ə�ky�����7�2�p��d���("-��M�Py��t��@L�my��6|�=