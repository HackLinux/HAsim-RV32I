>�<��3M�"b{�t�̶'Y��k��M��n�}�`^J㒩�CU�ޒˇ��2�pO��ʀ8|�5��j��FE��!��>D�1C%�8p�9V��?��#e��t��&����D����d��֕��Rd�8�7u�L���+mߕs��� bz�C��0�U���R!�&Ô%c�!9ۼ	�4��˵�p��T����A���;B��I�������T��;��|���;m�k���)x���|�}��d���Tl�;�S�����$0��,�	R�
����`�A�^b�_��\U�$$�Z�o��_��)��uz����S9�$�]�Ըْ>�Ћ����$�U�ʆ��U�W2��A��f�z&��:@������UV�N�0�w<E�i?P�l�y��e�8v�։�`����N�7��n���d��3~�5F,$Ag�^gQ�c��iSi����R_�E�J�9䔑�%-w&�#b��[�Q0���6�9)S�`�Tl�W&'7���*��Q�QS�����]T��9������P�d�� s�c���X
k�R:�p#Ƞ����J��(��O���4T�$B]u��z
�֍�dE�W�,����"�As.��XŎYs�s��y��dD�3��[B1_'��>z �R�y�$�l�M�&9�7Qa�d�^�?{	��A[��T��hW1�;1� ���h��م����r�c0P��6�$�<�����"�㶮܎2�Aý�<���~�#��;��÷�{։�J"�xE��S	b�~�bg���,�{���~�i�ق9�8��|D�Q<��?�IxΏ5 �j�����+�:ԫ2��CO >�0,~UҏC�;z��&\���;��?��^b)ي#4$�*�����ӆ8���<�
�+R?�%�]���@���~,U[�e`�oa�$�3� ���1CaD�T�-oH�u�O�o���~���I�hb�O��L/��Q�u["�qǎ����~�\�قK���5�z�4J��%��2�)y��!�$��;��)�oͻ��j1�vB��BÏ9{�X�i�� gcm��8�_���Ҍ-?|�kb�i�����|�E0XJrQը5�X/��+�sFs�#e��lS�I������4��<~�(��}��gZ��Ќ�f���[��e��o�n�Z�&7�;�˗��X�� P�B�3p۲S�[����e��6b�VR碩7�&(P��.�X:���Y��|> �v��� &��
�=�!]�*����R�Ķ%�)��j�%Z��_�Q�m�����X�����~�^�_�?�e}��c���{��-W,E����埠A�2�O�� R����D�i(��P|'���
��1�aMo,|;�Gl�y'R����\������h'���T/��?�cBڪ�#b�vI�E$�?din�r}����W8��������H�kK�]�-M�e�4�&Z��c�i�3�V��R�h�+������>]c� �e�@�L[B���/�6<�$�/��T�%O\q��w�E����{��3��o��o��<6N�䂾�<�9��:ժ��h�lۢ��I�畟��%�Oc���5��YŎYs���8(P�h����$>S�3P��A�3�7�c�&������f�1����Z�b����5�7�E��"v���܄�n֮��:ܓ<6�=��F�