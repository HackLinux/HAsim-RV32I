������|=J�������������������+v�������������������ov�������������������������ߎk}n���������������������� �Y� ����������������� /5��������������������}������������������� t(������������������� .������������������� �fc��������������������#�\������������������p��������������������3#g������������������ �������������������������}��T�|j}��������������������� �[V ������������������w��������������������p���������������������bEV������������������� �â������������������ �%��������������������#Ng������������������W$�������������������L�g�������������������d�c������������������������꿒*9O��������������������� ��� ����������������� �E���������������������V ������������������ ���������������������� ��������������������� ����������������������2�#K������������������mF������������������� 4����������������������K��������������������L���j)���������������������� �:��������������������կ���������������������抢������������������������������������������)6s������������������ ݋��������������������"0cg������������������59��������������������f��������������������� �K��������������������/�����jRR������������������������J!!������������������������������������������#���������������������4i��������������������f������������������� �����������������������3vf�������������������f3���������������������K��������������������ԇ����������������������*���kjk���������������������� �4#����������������� ��x������������������� �K%������������������ L0c;���������������������d������������������ $!!��������������������4J�������������������h�f���������������������0������������������ �����������������������ܽ�� �@*97����������������������޴��������������������޽���������������������Բ�������������������޽�����������������������������������������������������������������������ƣ���������������޽����������������������製�������������������޽������������������Ɨ���b �np5(��ŎɎ���펿�������Ш��Ш��٨���𩮧�m����T�mm�������R}��٭�٩��������٦ѭ��y(�99mw�w�m�O�����OOQ>||@}�����V�>�})OOOQ>@@�n+*+ѭk�jUnQ�jnn*�*n�En+U,�j��XnU�nUn�j�j||U+�j::n:�pU���:�nn:U�|��pn̯n��������n��������|RR��e���h�����O���d��}������*I*���с��n�����ҝ+@G]_],,p�_����}��^G�CDUC,WWC�pC..,,pW�pW�U����Zq�������Wp.YX.W,,X���W�W�UWD�DYX�XX�.X+AB@*+����>+)��}++R@)|U�U|��n@nn�*p++�U�*>99On<n*���|h�()|ROpj����U=��������nW����nU�����p�U=::46v�v O�������"m5�b���׽�t��ݴ��I`HI1��((e7(utuX�e(��շ��e�L466JL64JJ075(77��yh���Le4�e�O��e����𬬷���L�dPJ3d/!33�666<'! 3��hO6J)8O�����e����a74J344hhh)ea")O9(>�7�V�O@R}}���()�m�V}>|eL(m97e4L�Oy��4J32�|3�������|>)aaa/2 s��Ͳ���v@R)�}}�*�}R}-R��-EEEC��E���E��E^�.^F^�C^F,W���^.G^GGG��G_��D����]]___]Y]]Dq�]_]DXXW�DY�YqYDXXXDDYDq�YZ�XXXXWXA�A;i;=<'f��9)���������}>}�R�����}��@�}��}}}|���}�}*@j���@�}}>@������*�**@�}��@@*�@*@*|@}j|}9)Qjj@kk@|�QO��O�a�L33��e�t�QǒR����������
b�������R���
�
w����
����a�*ΒRh����������������������������������������<���������������������������������������f�������������������#�����������@�}9���������������������O���������&����������k���������a��������h��������������������f���������&����������f�����������k�|�����������mm�����������������������������n���������������������������������������P���������#����������d�������������|Re����������������������������������������k���������>��������9���������������������k���������#����������������������*�RRe���������w7��������E���������+��������������������7��������@���������������������8���������x����������f�����������*�>>a����������7��������*��������������������������������������������������������������z����������z����������#����������b�RR�����������(���������-���������U����������k����������}�������������������b����������p���������x��������������������w}��|a����������7��������U���������U����������*���������Q��������m����������w����������Mi���������z���������$O����������b*�|>5��������������������������������������������������)���������)�������������������������������4����������������������U�>|�9R}�����@ϑ�R})@���w�@�}>�}>�7�>R)}R>)()���e5hhh��>��6y6))9w7)e55aaae(eɦh344L�V6OMVhL66���j8�j4O�<�8�PP��6d44�0LJ�7�n�Q>����
�T������V�m5m��7��ǧ�����������|j����������m��������������������$,����������p��������|��������������������wQ��������������������:����������z����������5��R*�������������������������������W���������`���������}�������������������<��������������������z����������?�����������*M|k����������m��������T�����������A����������+��������)������������������w����������k����������=���������`:�����������*�|j�������������������������������������������������)��������������������Q���������~:���������tf����������:����������>�}j��������������������������������W�����������������������������m����������P����������i����������x���������`P�����������@�|���������������������������������B��������������������������)���������w<����������:����������:���������Č�����������}�@���������@���������b�����������W����������+��������O��������������������P����������:����������:����������P�����������k�}}��������������������������������.����������p���������Q��������������������P����������:���������`����������`?�����������j�}���������V���������������������X����������*��������@��������������������h����������p����������:����������=�����������}�@�9a�״5�b�b����"�u�5�5�ϩw7�757����979e�(7997�je(O)|�)7)`9mh�|R9(y(5wR��)e)�)�wbaeee�aL7Q$)Oh|)(�ɴ$O��2�/�u���L�����eaa��쒠���>���>)+U*(��kk>)n��-��*n@|yRR��p@||}|n*�5+�R|>@}��I�@Q>(��kRn*++ne::��n��:**y�@Q@@@nn�U&�:x&&OQ�(:�dd6!����h�@�>+��
��
����D���
U�
m��k~�ܪ�:��`@@���������}���������������������Y����������p���������}��������m���������Ώ����������p����������{����������'����������wn`*����������������������������������������$p����������������9��������������������~p����������=����������z�����������+�������������������w�����������W����������.��������}���������V�����������Q����������p����������=���������`'����������5+�*U���������-���������������������X����������p��������k�������������������j���������wn����������<����������&����������w����������������������������������p����������p��������k�������������������=��������������������S����������=����������w��R����������������������������������������$,����������������R��������������������wn����������<����������:����������w+�*������������������������������wU����������W���������n��������|����������k����������+����������i����������<����������wU�>���������*���������������������p���������$C��������U���������������������Ϗ����������p���������`A����������i����������wn�*>����������b�������������������@���������n��������>��������V�������������������w����������M�����������������������n`���|��(|>@R�(>>OQ<jw9Cn>|U����k>n�*-�Rɓ*�n���*��QUnnnUU�CV��}+nUCU,nw+n+�+}+U�)�**nnUP��w�f8f8d8O8PaOLL4L6v4J��w��@��eLe(��e�ח��eaua5a�ؗmm557�7�����@�a7e���w��+w7���7���T@5�(�e�7bb��9�a75������ube�5"��4wh�((7��ӽ�nu/uss�IIu����s��ɿӢ���`@�������������������������������������������C��������+������������������j���������wU���������`p����������;����������5U�*Q�������������������)����������wn������������������,������������������T����������U����������A����������=����������T�`nn���������E���������������������Q���������TU��������C�������������������>����������n����������n����������=����������T+�*����������}w���������R��������������������~W��������,����������������������������������������=����������������������U�*|���������7��������������������n������������������.������������������Tj����������n���������`�����������n����������U�n���������-�����������������������������wC��������W�������������������n���������������������A���������`������������U�n|���������-���������9�����������k����������n���������,��������p���������wn�������������������`A����������P����������wU��U����������T���������������������|����������U��������U�������������������k���������wn����������S����������x����������wj�*+�������������������|���������������������΀���������@��������������������Q����������n����������?����������'�����������n�n�����
���w��p�������������±����±�j�����±�b�������}���±����`3�n�*-�5�7����5���m��5��577�w�57����7�5b��777�w55���w5���75����w�؉75����5�5��55�����״�5���5�5�ʉ��57�5�5��5ea777797��"7555�5u"a�}�*}���������+���������9����������mV���������π��������,��������n���������7R����������}���������M?����������&�����������*�-���������pb������������������m����������w�����������������������������<���������ئ���������ߏ����������x������������$k����������C����������O����������>���������b���������?��������n��������������������������������?����������&�����������p�}U����������nb��������>��������������������U���������W��������C�����������n����������=����������?����������P�������������>*������������������O��������������������+���������p��������U���������m>����������n����������i����������P�����������U�}+���������U���������9���������������������U��������U��������+����������>���������،����������z����������k����������mU�}*���������*���������)���������w)����������U��������U��������U����������V6���������7z������������������~P����������(+�|����������n�������������������w����������������������������W���������@���������������������=����������O�����������n�}k���������U~��������O����������V����������U��������*��������U����������m(����������h����������A���������~�����������9��|�����������-���������R���������7�����������U���������+���������*���������������������+���������~:���������~:�������������}m7m�9���7(�)�4LLhee��yR@}RR>}|55�>)>>|}|)�U�}9>j}>*��j��Q<R@n+��k�}>n@k>w�+|j>8��|>R>j@RQQj$��888�O�Q��L26y93L"��5��}�����au���bꮿt1I1HI"��)wub5�I5wƥɩ55��׈����*w5��7�7ؿ�4���e�e���Ŏ�"����μ���7��"Itt$t6�k47�e�"�ŽM4�����u����a�uޅ�/��`ɗ��j|���������E���������P���������m�����������W��������U���������U����������7����������8���������:���������T�����������y��|j����������~��������j���������yV����������U����������������k����������m����������w���������TQ����������4�������������}���������*~��������@���������������������U��������p��������n���������)����������R���������w�����������4����������yU�O��������������������}�����������������������������W��������k����������)1����������n����������v���������be�������������@���������������������������VV���������$C�������������������������b�����������Q����������6���������������������y��k���������@~�����������������������������j���������*�����������������h"��������������������4����������a����������j��j����������V~��������O�����������������������������n��������>����������>a����������6��������������������9a����������Q�|Q���������������������������m����������$*�����������������h���������l����������>����������&���������������������4}�)���������������������)�����������������������������)������������������2c����������m��������������������I�����������J�})����������#��������������������K�������������������d������������������J3����������v���������·������������������������n7�ݴw�Ɨ�w������׈�����w�؈�7���7���؊�e5�5�ɿ�ؾ����7�ب����e�7�9���(���h�(�yy��})y9h�7(��yh�yyh�yh����hy��������e��a�Չ����ʅn7�V���ѩ�(7@|��}���k>j:|kjQP�U�>**nn�k���k�n}kU��nP<Q=6�QQhQ|}Ryy>OQ�@jQ�||@V�eO@�}�)�)RjP�>QQ��RQjk�Q�Qj4LLaa�͇|(|@@|�|�@--**nn+EE+UU�UUC�C�pppCCE,,pp�U?pppCp===kPf&&64�|��������������e�������������w����)���������V���������(�����������������������������������������V��������7�������������������������(��������������m������������������������������������������������Q���������������������(���������������������������������|���V�m�VV�RVV��5��7��9��V����7m��m������(����5w��j�����m�������������9��������������(���������e���������7j������������������9���������V����9����������������������������������(������������h������������������7@�����m�������������9����V���������O���������e���������������������������5�@V���>VV����ڊ���Бm�m���@)�m큩}�O�}V��n��mV�>RO�mO77�77��������������������9���������������(������������������n�����������������>�����������������������h��������(}���������}����������)���������������h����������h�����������|�������������������V��������������9���������9������������V��9��@�����±(��������*>��9�>m(���k�����������������������-����V�������������������������9k����m��������������9����������������9���������h���������7k�����������>������������������������)���������h��������9n��������������������������������)���������9�������