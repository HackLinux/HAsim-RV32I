v����pA=Sm����������eHLTw�Ϊh45\{��������~tpLGry{��������f\ORl����}Qf�w�����w��h~�TRkj�����{���|VNZf�����8Tzy�����u�mpZ;F[y���������lRKPi����c/Upq��������~�iG`ky��������~q^bq|��ʶ`Jng����y��ow�\IY{�����pws{�gYW_���Ȏ1=gk�����z��vvhFBb�����zx����ogjw����d1Mfc�����w���v\FYn}����|����~nkt����O>^f�«��y��|}S>^�����|p{���zmjk����y3Ht������|���mF)5h�����s����yh`ep���nC3Qn����y~����uC?w������~���{}rpx~���_=[mp����s{����e<Oy�����in�}uufepu���mEES��Ħ�lg����e,:Y��̷�oY}��rrnx����u3Zh�̨�yaw����A)c��ñ�tcg��se_`�����+Mi�Ⱦ��rp����_6T�����jm���r^r�����Q:hz�ɤ��s����yJWn{����tgu���sfq����a-9NS��ĕ�{�����TAb�����c`ox��hXe}����H-;x�����x��|�d.6Rz����l^o����YN����oB[�Ὺ�q���wo6%d������_a����oYu���j)7_��آ�����rnN)K������li����wip���y0+V�����xx���tK;e��Ż�w^ey��rqy����M0DOg�Ʈ�`k���wJ?Nb��Ա�Wb{{��spz����K*7i�ͤ�q[����`9[���pWQf����kn����\%+W�⹝{[l��~?#*Z���ЋW^w���vhm����#+_��Ȝ�uo|��m8"C���®�jg����wo����^>Br�Ĳ��iu���S6H[���ӎPWn���pgc|���@'09�յ�e[s{��b<K���Ͷva}���}Y`h���W)U��̻�az����31Da��Ժ�lds{�}_Xw��ٛ3r�ʤ�|ntw��m2Hcy��Ȭz^qy}��af~���Y(K��Ʋ�]k����QMaa��˿�^c����obp��ũ9	_�ױ�l_�{��}>HYn�˺�uls���{i`���Ҏ&6R��ȸ�z{����Z;Jdx����yr��{qkn{���`*'"9�ؾ��oy�}��KHUU�����qt����xnr{���],8/[���đt}o��}=EXf������|��x{yssr���`5-*O�����|c^|�yPNbgr����wz�|��~ymg�ɿ�h2'f��ؽ�uie��vTNZfr�����}tpm}�yol}���E 5b�Ű�{QXgp�Ygja��ƹ�vlv����nr|���` $X��Կ�gd`r��VRah������slo���puz���k)&Cz�ǲ�G?m��xhkkq�����ssu����ys����c!)<`�־��bTZs�wjfn�������ibiq�z�����r@.AVo�˽�YIFXw}~|�������u]gqw��|�����SAAZ}�����iMU\o��z�������RW\i�����~���jWWVs����eOTTi������|����o][j}����xu��z`\df|����rRKUv���~xm��}`_^h�����z���y[NHZ����zgXd����}t|����{r`d�����qt���xXQWc����kSIm����zt�����}r^d~����pw����;4MY�����bUfv�����wx����t^fv����rsx���MKNN�Ĺ��WLRh����|x}vy��xko�����oyq��x3/6N�����hXTj�����}�z{����xy�����}w���^DVlw�¹�wZMl����suuel���|w���xzuv���m5;jv���sddbg}���{ywmk|����������wy���]8R|����k_[`����sxrmt����~������wn��vI9To~���a[Xc{���}ovpqx���������������gDK����s`]gx����wnpqlv���{������}�lL?=Y�����hgku{����klku}���{{���������lUUe~����wjty�����|hjjpy���|}y����kcc^P\v��||x������yquy����~v�����pktrlw��|rr�����������wnhn{���~iu����}l_aox}�x`a~����yww���~ui`z����rm}����jdfp����ir���~|�����xsnev��|ndv����wjis{y|��nhs|����zuy���vpqrz���t{������xv�����sv����~��~���|qsxt���qor����zjer{�qcfs������~�����oix|���knvy�����|~����qq�����oy������veems|}rorm}���wnkuxx|n^m����|{~{���{z|p}��tgi|������zy����ziiy����|wy�����zlj��khsy{����pfhoy~uij����}nt~���~mr{���tiir������x����tv{����pz�����mt�r]`cp������ymnzujkns����}~���~~��~ukkpu���������~}tn{������������yx���pddein���{����uuj`oxt��|xy~��yyzxy���hbnut�����������mbk������{����xtyw���wRYco����rp����y[UZ`{���{oo|���vqss���f\jko����{�����}hhpu�����y�����msy}���ue^_i���ylw����~dVViy���zrxx{�zstt|���mkjl�����|�����qhhis|�����{}{}������rmjn~���������wc_abfq���}xwstuu|������wnifv����������tnrqpz�����wrpw�������{uvlm{���������pb`fbao}���zsmiqx~������qoki}���������~prwpr�����ymknw�������idhgt���������vgeilji~���tqmkt}�������tjnml��������zwtuz{�����}{vsv�������iefgm|�������{qomhnqq���wqttt|�������zvsnj�������|ovyuyy~���}}�vmii~��������xgk�������yspomjv����xsvxqkr�������y��|iq��������tstv~������~��xpnr�����zx���nn~~z����zqignx����|pr|xsonv�����x}����mv��������vmm�����}x}yvsnw��yqy���tr{{v�����vkchz�����zrrrsw|���uv~����~|����~�����~lp|�����ypouyx}��~mnz����{s��vwvw����vgmtz����ykjhp~���wmy�����zu���y�����~ws{�����uppnqx���zuv~���u~���rt����xqenxy����uddhq���ysr|����wt���|�������}|�~����{yriem|��{wwx{���u~��zqw���}zpsxu|���}vqfds���}z������y���y������w{{z�����rkcf|��yqmz���|v���ww}���yrpz||���{trgdiu|�|w~������}��}is������sr�������xtmgu��|tpv����~tw��zr{����~{uvz}�����urkj}��yqit�����z|���������}}������wngr��xjiq{���~tw��vu{���{|}xw}������{kdr���~ml�����yu���}����r{�}��������|wtpqsxytt{������}��}}���zvw|}}�������|kffj{�ytpr����wt}�������~~�����������|lhtzzurtz~�����|{|����rmpv����������ueblsvxyz{|��������{�����xvyz��������ywogkstonw����}v|�{q~����sqw~������ztnhiinutw������ww���~������~mk�������uopnorupkjw�����rs~��~~���|yzyuw}�����njjddnz�ymy����wis���������|xuz������|ohihn|yqu������qjz���~����{utx}�����{j``gq�|y�����{qp~��������{smo|�����}ssnhjr�{mu�����vns���~}���qgbdz�����~rmi`bv��|}�����{kk���������pdo��������|vmdgm|�zz������wx��}vx���vibjy�������|r`Wew��|����yjr���}����ycdj��������tpmflx~�wq|����thx��������qhfm{������vnkfggt�~{������sk���������xnp��������ujglu~�yks����~kkt|������}mllv�������korg\_p{wv�����wju���������}sstz������ysojeiwztx�����uks��������ypnx�������xtoaXanrqz�����vlq��������ztrs��������z|n_[izskx�����wqx��������{sqqp~������zncZZnwqsx�����mt��������~qry��������|tcPWirwtt����{mcn~{�����xsmq{��������q^S`svp{������tk{��}�����wqtw��������zpe\cosvt{�����ifu�|u�����uqnq|������zkWZdmvmdv�����sz��������ztrqs��������|f[_kmdfp|�����nv��������{sqms�������tnm^\\Y_el������v�������~txwsx�������ushZNN[ap�������{��}wz��}}~{uq������qk]GDMZr�������������y������~�������ja_SFKi����������puwpy������~{{�����`PUXZU^w���������{kp~��������tz����tomhq|k[i{��������wjev��������ysk~�yefpomuze\m����������}}���������~|rfk{wr���|yoci���|ts�����|y���������aJN`n����txylinqvro~�����}��������_SUW`u���������lX_v}��������yzz��z\Zgggwuoz������v[Z[Yj����������wr�eTYfv���{vw������uefmpr{����������SFXbm|����}�����v|�|vtuqeh��������eUOQc����������tly������wwzts|����jNftt}xu��x�����qlmfp��������~jbgpkRATgt�����u����|{��y�������������|<%FWl����������vYbks��������������P1486In���������l[irx��������������`Z`Vcvk\gx������v��qmt��|�������{CCZ_j���umg_e{�|hjw����u{��������r?CSY}������}v~mWnyr��������}������uW__cwx��������PFQNfy��������xp��oFZtv��|z}z�����zobW]`hu�����������NC_[f�����~����hfwzzxnhYRi���������ZHEC]����������eg~������jkjq�������Mc{jv~t��������[]h`q������{xo]Xd�k?Q`b�����x��������ow}~��������kv�e28V[c������x��teq�����{wu���������g:-5V����������uUht|�����{}z�������{C7B8;f���������|g^]y���������us����]GP<5Tdhv��������|rei����������yv��}GRf\fzxzyr����p{�����y������������oGNSDj��trhgs���|mt�����ml���������_<JPT�����ux|��wfrxw�����xwx��������R369N�������zxpKImsv���������zl|����`HKA]���������qPFOYp���������w`q����HTl^s����������LISMZk~��������zpt���iGW|�����{�����hac`qxp|�������������J>RGpĿ��to����zo|sqzzq[^�����x����z<>PM{�������{��uo����uibfo���������c>ADS���������bh|v����r]bhgy�w}����eOG9L����������\Wq|�����fijirgi�����fEOX`t���������u\idn�����}vhi_Nd����\>V_r��gm�������jxy~�������}fWfx���d@IPh���qdr����~j~��~hpz����|f[cx��mG@Sh�����~����fp����yqhw�����xw|��wA=W]|�������tzyYSu����~tt}���~|����r0 5Q{���������uWVp~�������x��vs����r""Kj���������yN>Rj}�������zsvqp{���x5Bo���������|DAf����������vjjv�����42Uc����������\Qbhq���������_Y�����ABSPu�rv������~MXojv���������~so�����FWld��xmx�����gYmu{�~}~y������x�����:9`j}�rdic�����^_rn���{zy�����������G<N^y���ts�����k_vzy��~xpv�����������.%DMw��zxsz~n��dWq|���vwv���������ɓF#+En���������zf\m���qu|�����tr���Α(BMx��~�����oY<Kqz���lh�����{z���ȗP5BRh���������zUA_|����������zon�����@9`ew�tx�����}V49Rh~���������tgn����OOsm��wav}����xFDis}���������~xw����|F[z}��yjn{���uRSsupxvz������xag����}:Mlz�����nz|y�~exv��}�������rw����i<M_r����yxgc}tew���ywqr�����w�����QBZ_}�������~wob{�����}�������}�����PCZXm��k}�����|PUx����|���lqox����wILULh�yt�������jnnaw�������xshr����i7GSZv|kp������dgufbr�������qp|���L->D\�{ruu�����}g~��xm{�������x����WJ\b{��{�������Og����wqlk�����y����O&>^i}ip������ri~����������������{BAZR^��tt������[a����{������pkp���z40^[a{ih�������WZzu~����������}����dJio}��cpz�����vm��{�|o�����������f4Cli��nx����}�yQm��{lp������������a2Wb��������|jJY��y{}����~y������`BKPNYeeo������cWmpq}ut���������À)8opw�kdty�����ko�mnmm������������{0>ZMt�vdy������|����pct{����������A'2If��~�������a_y��������~u{������TMPF^ubn�������v�y^eim������������x6P`I\h]y����������mhZa~����������P BtlomFM�������q���}\]u{��p�������[ 8BS�}Wg������]q����p{�����������wNUUPc`OZo������y��|{x�����������W]}tonXe�}v��������skgv�����������4,NYp�ii�����zpg���|v����}m������dLX_\]\TVx�����pdiq|�wu�������z���t7Poivwbhtx�����|�~eefu�����������`@JZ[cfYe����x�����zqkl��}~������xLC\`cs^Os������}����ss�����vy�����:,Lanxk^i������it��~ljw����������xD=PTeqZYr������������������������|1)JPXb`g������qz��x{�����plx������UI\M@POMs������ql~�|||������������TNhddlPJk������t�qpnt�������������TOuxpo]Wcn~����oy��y{vz������������aEUdkunj{���op~tx�yq|��������������`V]STbip������n[Zoxko~�����~t�������r`wjftir������ckzij|������}��������bZgWYrf_{������y}[]sz�������������sOXh]fur|���������|mmkt�������������^EOVV`iny�����wt��}rptu{�����������X:9BWjpv������b[�����wy~|{��������i9+;Wiszz������fT]q������}vtr}�������B,;6Ipxw������}ihqox�������stvs�����c=8DRYk}}������nanvde������{mifh�����F1O^^f_^}�����zjm|~wu}�����|rfi{����vL7Qfds|jo�����zn~��}yx�����winqx����rHOdW`qgfp������u������}����������~�mF]jVl�wz������~���|�����|}������}ht|WPo_Gdvoy������|��������{}������y�|KNi^f�rc������������|��~x��������gCM[Qgzeq����mrns��������������������qMON\�~cr������io�������������}������M>TKTym^r������\j������������so�����^;YaXigRf������}x}t{���������sio~����_\^NRWDW����������pv����������������s{rXWVC@a�����}�����lf�������������qVfro_E@Oe�����z������}u������������QNe_h|iT]gy�������|v�����ghx��������W\aSXbk~�|�����~��ru�����ke��������zvbKIMTo���������{}�����x{�~�����ttuZGSQCPs������w~vnz����tz���������s�ziqdSdt~�������it~�~v{zs~������ZcycYd\_qw�����x�������zmqm{�������dw~VPabs���������t|����qls������rVmyb[[NGVw��������{rt���{���������umxiYc_Oa��x�������rw��|gbn~������odqfZ\XOau��������x|���ynil�������{xbRB:Mjy�������dg����{w{�������g���][VTglv��������|�|z�zw}�������n\lschtljvxzuv�����r����|ROq����������eKXTd�������z~��tx��}nryvw������p}xcicDFm��������fk���unno��������i{}gtvdork}�������qw�vmw|t}�������wiwn\eo`^t����������tkajvfUr��������mQSY_bel�������y�������|}zpp�������o`pbDEVai}���������aVu����is��|�����zSevcYRW{���������}NSes�������������l?[g^pgDS����������y`Uj~�������������nYj_Xkfe�������z��s~w}������������mOdlX_b[p�����um���uow��yz{���������h\tiam`i����{~�s���qz����yjx��������~.5f`_se^���mf|~{��}}����uTg���������9 Xol}s[m���rv�|n���������oZq��������a/@nlhw]H���}tqy����������ol}���������XHceizkcw���tv}|���������uu���������v/Dc^dh]`z��~ry����yz�����qs���������Z6HQVb_chs����ws��tsx�����yr����������M>GKWfWR{����ocl�t}������zz���������cDIJQkg\{����|jr��~v�������}~��|�����g-DNJ```{�����wiw��ot������zu{yz����|*0PNR\NW������wgo��ti�����|ry{w~�����0+^YEQVUt���wzwrx��}|����}}��|x����d/2MMK\^Ro���}~�wp~}y����������t����A'XiRPNJZ������yxtq������}���~}���a26QTPWVUp��������snl����������������K9OKI\VLg��z�����d\m���������������OC^\EBMRc��ws�����oZ}��x�����������i_u^EH7=n���x�������sw�~o�������Į{ez�kNF>Gr�vs����������gips��������{e��dKRE:f�p_����������zR\ir��������eeo]FKRN\ql^]t��|�������skww}tl���ŗ{�y9@QTr~y]g�row�������tjrcerz�ђ|���W59g��}uw��eo{��������odv�����u}��uX:Ei~�xl}��sgip��~����xjs���fF���]pqipvz����x~~zwwxvpx���������I_��kdfr��x\m����������gg{wlm{�����RMmbRUNQv��g\���������sen~~ysr�����u~��ZIYit��������������\T^q�{qt����cBn�mAGVktknr���������^_mms}�����xT[urVBQw�{bj����z������wkv{xsl~����pl�d7?H`~��z]|��r[�����|p��{pj�����}��W?EFNl������{v�����v}��nct�����hf||H-GKEi�������gy��������ifo�����MF��E+6FTt��������~v��������ru}�����JX��?+@[^h���������yi}��zpz�wlv�����QY�|B2=Ww~~��������}t������}}qp����}[}}G:APo���������~xz��z����l[j}����Cg�vEO^am����������zz���}���sekl�����cu�[Rabkqx��������xz������wsmied~���jw�~PUddju������sw}�����~wolqoo�����nu�`KU]bt���q���vz�������{|oimoz������uxnaVOc���{p���thx����{q}|mdccx�����{m��hXYj���������s}����~���xji������wk��dJT]q��z���zfr�~snqpopk\Wfz������u]erXGTYVj���~{��}��l|����������������m����|x������������rt�}v~�xu}��������QEioH7GKYswmhgdR:DTA0F]`ec]ev��r}�����l���������ű������}|����������������Ücp��nfcn���}xupbI89BLY]SMV]Xae\_p����}_t�yW^g�������|j`pyj���s��������˶����z��o~������u��\DJScz�q_hwh]jqnow����oK_wbFJdw~�r_r�yPRfkhp��zl������������������xtv���������ks~���{�������z�����GC_R@:@\s~�qdstqo]\`a��vz����uu��������aZwaHU[|���}���|ml��������������������qKLR>Kj^QcqsnlwvcZ^q}u}�}|��������z}���hG>c{eY`^j���������}y�������������������G6]`C@PXm��vvywvl^`mx����}|���{x��������<8gun_Qa����yw���uv����������������������MPVJ]oip��ykglrk\aicp�s{�}{���~~������rRu�lv~no���xx��{ylku���w����������������]_r\PW\cq��tiquwvg_k}���~|��yhjp��������YG[a[^Z[clz��yy���~rey��y~���������������m]kmSSkeh������yuti^p���~~���spty���z|x^HZsmkrqu���sQY���zttw���x������rfx����ĩ�����y{��������qjmr}zt|���{ldbkx~������RU|xiomn{���qeuynidc���phcw����z��������~����{w����spxpnuaQcz~tgr����{�|||�����R?q�oje^s���uq}���bUQo��w}����������������hT~����u}���{v{yphb]e{��~�����dQ_q}�����}QEl|_Up����}qy��z|�������xwxw��~����������hn���}vdr��������y^GRmslc_k���y{�~v���t��sFUol~�uh����xny�{tij{����������ynq������Ò?Hw{{�������{tmjs|vcd}��~wsy�������}lgh}��JAs~gaedo����ux��qo{���������|\h��xw�����pDHk��zm{����}�����~v{��seXVfks{ncfkxla����p6evGRjay����||����hS^y��yu����������������u_�����������v��wmqjbkw~{u�����{uyuvwr}����GS�lMU`kvrz}dW_emnioz���}������yw|}�������sWk���j]w�������������~���������~||~ig����e&AhYGPf~����pswux^GQgr~�ws����ztuz����t���|q�����������������ysx����y����zd`o{}�����ZMd^HU_Zdq��sgqkjysqyic�����zw������������jc��v���������������}�������pntqiku|}}��i"8f]\j`h����vq|��tVWai{�v}����wor����x����u�����o���õ�x�z��gg{��������smow|�������d*O~mbbICb���|~tlroh\\n}}}�����xr�����|���G?np\flv������������������������xx�����~��WKy|cbW\y��������zb\\m��t~�|pq~}piighny���sV����x���¤���������������}snnt{vv�����[Nnup�|\Vk���~}zsmi`evtgnumdu���zv��������Li�vgu{���������vtzp\q������������������yEP��kj\Xs����elrl`QWo~����������|xvus|����lVju�war����������������������zuqu������em�cP\]gy���~��y{uk_dsiVdunivz}�~{�����qL\uoknqw|��������gfnls�����������������{Hg�xljYl����}{w\Vfi_Xh�������}spa]luz����jCd�j`k]`���������y�������������zz�������mMs�tszin���yx�wwria_t�zuxsvypgimssx����|SPq}puy|�������t|�vms����������z{�������uo�}aafdo����w��xvl\`l�����~z}�|tz������h7X{okxpoz������wn|�res��|�������y~������sV^wwjv}qt���|���txtks���������u`k{������bl�p_f`[s����s�~��dSh���wvu���vu��������ie��w�yo{�����}rvth^e~���������s~������}H\�ym}zomr��wmrgg��se{�����������~yw�����WUokW]kfe|������p|��uq��������}ov~�����iGSgUM`hs��������uyzu������������y������k^��{srg�����s���tnnqy��������xspnu||���p3O�ughW_���|k~�pftraaw�s������}~�������rf|~lmss|����o��sr]G`����������n^go}����Zbi\XYT]u����qkjgz�rz����������h`jy������m��{hg_x��������chear�����������ymbco|��p=Jvvilfl����rp�iilVGo����������}txsq����aSu�{vxmy���������g`b`r�z|����}�����x����|RIef^jow����zz�{mqWBNepsw{��������������vXQbifqpn��������|��ee�����������rv������|aR_YARj`h�������nw}n`Zfw{}����|�������rBIcVL[jx�����������}vs|��yw{���xrx�������\LZWXkd_��������usumhmohhkebkt������������RQg^T\X^v��������}kd\d��|�����������������iSht^WXJV���yv��~}�}jcs|g_puqw~y|���������[7VeUSW[`i�����������t}��x���������������vIUh]bbNSgr���������oct�{ocbjmpmfp���������lcppfkjer�����������or~|th_r��������������pZ^[W\]Z\by�}pysiy�~rs��|]Nq���{my���������lvwikgY[j����������������ms��uj{��������cALdVVgb_m{�����������~�}ofag{��slny������kmyeakltz���������������zhVh��|~{��������u]u�qgcV_~�uhfpqoppnrw����wb^ijt|rr��������wu�zehna\aqwnfr������������}|��|z��������vOKWZTYc_cw���urw���~�����r]huvshejr{|������Wi~wj\^svs}zw������������odmtocl����������n��tfov{�nr}��}y�����wklnhfeefr��������udmrmaQUgnql^`ef{��{����~x~�����~���������SPkd`aU`s|�xzut��|�������}zux{}~��������u\y�thZHWx�rbdilx�����������{uroqt~��������ae�usfius��wmrit���������~zupz�~z��������zhyywbR`pz~oddUVt�����������w������������bk}ooua[k~�owp[m���{������|��������}����zeo~yz|pjo|�}_giYh��xx����������}}vu{�����od~zq~vlmr��hqpXeupojn������������{r|�����br��s��z~{��siuog^UZgy�������������������jMq~qyumrv��ibmkeYSZ]j�����������wwrq�|�ySh�|��}�����uodOKPNH^����������y{�yx����pQp�}�hm���sm|fM]lhRMs�������������y����uWYidbu��������va\YJ?C[x������������������[Z|~sm`at����vefiSGMKWz��|��������������r?Uu^ZgZh�������gv�c>8Kc`_{��������������}N=Xhb`p|~�����q{x_I>Jfpr}~����{|�������yo�x`]\Zq�������uvu[BBYptsos��������������Nd�j]bNUs����}�twwcXTYigeogp���������ú�UVa\\fg]b���sy����qmq}|tndz����z��������on�kWbbV^x����{v��jbs����}q��wi��������Xjpd_bpww��vwxv��{z�������wzunmmqv�����nh�u[dis�����{vhiwrf`x�����}xqhb^ahg|����yc~�}vvdo������~Xfwhew��������t]WYWi������w���sk`x�������ehyi`eo��������c]VS^m�����bk��}�nl������nd[IIRh���������jZ\`Zk����rYo|��vw������xhbXQ\y����������ncefjn����{��{w��w�������sqnXPW`r���������~ichlir�PZ�zaijlpm�����zqoZQVi��������������������kz�������������ynjbcfruv�������~�o\agX[p_08_e_[R]b`ihbl_SVG9?CYqx������������������qv����������������ztpz�������������tpsvstf>7`mjpbZinspeps\[^OJAHckjzoft|{�~��sjswt|~aTu�����������������y��������������wrzuo�\a���|jktqvyx�{`WUNLMMYfs}|uqqwwxnSTa]cmqkRRx��}�������������z���������ƾ�����}vx����]x����vmki|���zhnhQIFTs|��r��~k]UNSRQd|~hSayh]kj_\l�����u~�rir��������ͻ�����~|�������{}�mW\{��|�|szsa^em���������vqU>HOPbos~yh_ea]ZP=;Y��|uvgcsphs~����ǿ�������up~������{����yQRz������y~zor{���������bVURLQh~���zZSZVL:1:Jc}{ha^VZaai~�����������tum[p�����Қt��ohacq{�������������������|sc^]MNrz�����WEO?6CLRc}��kgeKA^~�~��������|vrk_^v�����ӹ�klnjx���������tr�����������tehl`V`lw������83OLUicX^bde[URNaz}mj|����wdgkg_`rvy��������Vfy{���������������������uabpsns�{v�������a:Wtfhtfcj`adfw}pr{z~yv���u]^n`PWcgi{�������q}�y~�{}�z����������������ruypt~~���������vRdpYZZJMLRjem�~Wn��ueo}{uc`cZ[hiem�������P?`hftj\co��������°�������u���������������j_�zmqRF_o~~p~l���sh`q��uWMZ]^d`^hz�����|CDfc_`G?Ib��w��v�����������u{�������������q}zn{oXTXkugpyo������|z�}gV\``]epfc������fSYP>BIA<Kblfjqis�������~��ugz�����������ĕ���t~��wx�����vw���������xiaea[hu|�������on}eNRJFPX_b^prZ`urrz���|{tgchdbimw�����࿕�����xr���u��������������sukdcbfgh������~��rvkLE[nkRMYSS`^Zcw�����u^]^[WKDUeq�����������������������������Ͽ���{txrifs����|`h���zvt~lcebb_]ZRNamw�����yu[@CMPV^l�wZTjtmz�������wr�����r������������~wy������K]������������xYaki_OVglx��|��yodNIX`kv��S!9Q>Tzid������oiokbm��������������������ך_njZhiu���ž��ko}^LMUntmspr��vilics~~���hBGaQ>EDGk�������fVIOent����������������¨d^��uyt}����������qlosnr}���upvyk^n�����S6JI?PPKTe�mv�pes~yhiupmvsly������������ϰ�{�}js���������������������yu|�t\an���x���[8FJ>LVLRfwlOTldm��yeZn�ztlipv}xut{��������|�����������|�������������������vqvlkvx~���wS_topdROKUrpZWZ]jiegebhv�xhkrwztqhix������������~�|fn������|����������������yjdnqoru~����zV^^MPTIMg}g\RL]qlbcdip{xu|{olpibes������ͰhOfkiqtkr�����������}����ư�����mknt���������vRQbcedSO]u��mgfaidX_cl��p`holrofs��~vy}�����nUp{kjgdy��ū�z�����������wo������{yso}������^Mejehbk���lJTis��{qb]s�{tmw���~zqgjppy������xSv���sWQh���������}ys�������~ninywwz|{������[r�nIK]s���mj��qophbZr��rsu~ycbd`kldz��������c>Sxl_ikv����|����������x|���{u~�y���������GJt{rngx���fO]z����q]y��d][f~��zv�����uo{����^[}�|pjjs���������{kv�zlx��������vijnq|����{lq��pbal���~p����xZQi���zy���smvjjnisupz}�����yw�nUhw����p{���������rz��tjqvtx�{z~������br��mkwtrpfYc����������z_kvuvhcptnjes���������ku��`^`fy}{{����������gdtz}yhfkt�������������w�}^OUTXp�x����~}sl��rFPgpnbdrs|��{�y������`n��cfkr���t������ph���pz�������������������wo��|fesxri`bs��{cbgdt�yks}��vnmrkbl��lh�����aa����vu���p\aw����}w�ñ�����yvw��ln���x���������ve\g`WO?Hjxtnv�����ynlmpjdabicVS[euqq����q|��rm_Xn}vmeo����������������uptxgr���������kmjVOQLQdpjXc����}w��||{vqorsfVS\ddmy�������fRcvpiotw��������������������������������~{~t[QTblgk~���vyzsppxwq��y^l|zpq{|xxojk]OOUduvywkp����������w���������������������gfichnq�����v||{~{|�}|yppsqkhjmm}�����gei]VOFKV\bm~��������yw}���|mtv|�������������zst{yrpw�|mu�����v{��vtqrxvwzwroms{�����zbmxkb]cpuzqTRkno����������vt}�������{}���|������������|vpw��}���~������yt��}wrkaY\[\gv�|���zwvv~}pfs��w~������xy}}���x}���vh]as{x���������������xu~�{���pq���{vxxljkljkigbchnqq��w����yz}|zumnx���������{xz|sjkov��y���������������~���|~������zw}��zjcgjoqln{��{snqv������{w��~py��|twxojnwxx��yussy~}��������~������������|w{}{��~xy��~klsrquvy����������zeau�}u�������rhx�}lht~q^bopls~�������������}okkq}���~��sm|�zny��wimysfdq�������������yy��|vxwqx�~w{��{��zrnjfaX[lvplt���������~vx~�zsy�|xm`g}��������~nfjstqs~�������������yps|~ujhs��{vmi�����qay��so~��~}���������~{|xpjkkkornkt��|qnmw�vtwx~���w�����������������{qlnq~��z|���ybW]my{������������������ymq�s^folpvvrt{{trwwoifegp���������������qhgp~wiq������~��~}{rw}��}tz{y�������������zusj\S_t|yy��ymUMdp`Zent~��������������w���nddkmku��������xkdq��mn�����������������ow��{lr}}{vwwstsvyqbTS`ijkx����������}y{z�wkhm}������{miq|~~����wllv��������������k]aer}{vw���wrsxymdmyzvvzzqfn�������������uma\lzyy~��|fiw}}vw������������������~z}ytojdao��}~�|���vtx���tv��������vysntsx�������uuymhqxzuu}}rq}��}�������������spxkdmv~����}}wvsfhs~xjiuvsy����������������wjhe_fs}�������}|~wla[emq�������������{qw~~|uoliokdr���������~xtojdios}����{��������oknsusysjpqqvt����{y|vx}�����||����������wsvraX]mw{xrv|}rmotz���������������������x���pmroeft���~wy|sc\gsu}�������������������|}xy���u}�yllptqopla^ZYcq~��������������kcafqqipmez������xonpqxxtw{yy��������������~xsdVZeqwy�|x�����xxrbZblklqvwu{������������~zwspmcdmuw���s{���ts|whgt�������������������}���qhp|�����zv���pmurb]m���������y}�|{x{������~|}uos}���~m{���xs}�����������uoppossy����w���~tpou�{~�unw�zt}����}���ywpigditvvzzw���������|yuss{���}s�����������rowwsj`clklllu��������yuhcklm��������w|����pnqoppsod_ffnqq����������|tqv}���������}�sqx{qgmtutkjprtxy�����x����~ogkt}�������zupp��wjq{umlrw}wrwzx{�����������||us|���������tow|tgiy�uqx��|tvzxwz{���������|usoq{��������}mbjsnjm|��ux��ysvy{}}�����������tqt{��������{rmv�|~�}mix�{st|�}~|��������uqrkhjmt���~����wio|�~~���xw}�xnv��������������zywmhix��������|sq|}z����tu|rilmx��zq{��tv���~pllgksw���������lgx�}{��}vw��ypz���|uz������snuur~�����������||tgl�|yz}wlmuvw~xs����zstvut~��������������yutmjv��vouwvty}|{|{~���so��~������������������{rjbhqvzxv~|pc\frmv�������~u~������������������rdbt{rv{|m^gei{~z����w}�{{���������wqx�������}roy|tpw��zkfm����������������x��ztopx|�������i`gmnx����{rs|��������������|y|~~��}}�yq~�uzmjx������}sr~�������}��|���}��yr|�odv��x����yz~~����z{�������w{��}{����}j^ds}y����������z~����v{�xoqxwor������������uf_empy�|p���������|{~{rilwymb^`r��������}ws}�xmfbfswy�{y����������~zqmr|�tlns|�yq{��~wxp{��|q^]n|��������������gcnkhflw|vkgp~�~�����������sbau����|x�������~`hwvtvx���tq~��xu�����}����ztmgl|�~��fe�������wU]nnlnjw��yy��������������vhkot}��wot��������{`dwyqqy�����|��~��������n___^^co~�ytv~�����v]e{||������z�������zw��s\be\_kx��x{z~�������}qr{��������}u������}rpy��ttqghbd|�~y}���������yqlv������~yrr{����y��ur���qec`Vay}puzqn{���~��~vrv���yz��xw~������}}������~{����������������|����~}}��te{�wYQdtg_flrspjadtxuttvuqu{zyuobW^cY_u{ogt�tgottuvtogr�����������������������������������|{���jjjt{||}���uy|||s}�{iiomdgz~^FLU[leNWpn\QWe`Y``^^cny�����������������������������������wv�������������������pgjb[cnrsqwoRFSdhZSd_OUVS^iopfowkm�������|~|�ytz����������������������������������������||zonnghoz��z��ukmp_Q`qibgjbX[heYRYhf\ixvx}}vrwvkimlgiw���������������������������������������������ylx��x{zuvrmw��~ms��d]r�tbeoi_\bfiic]^bhlnx{bNbse[bnurqtz������������������������������������z���vv�����qr���z���d_swpijkd]]`djliglpigt{q`V_eYYa__gijju�v���up���~����|�������������������������������������{zyutstpdk��x^iy_EJWVPQX[]elmmw�sbv��nnxyfZbkibh�������������xtyvl{��������������������zttz~~������xfm~tUIWbXLV]]itspr||~��}ux|l\\[]b`][ithax��un��or��mjvv����������������������~|�������u��t����ppuqohj{���ihtppqr{zx}zsiYX_cd\S^np^Xkrc[gwvce|��zqu{|yq}���|��������������������������������������|y���tm|�racjpspiimrqs��oqvhYWUSSTfx{wrpq|�u`o���sv~tmfS\wxllw��������������������������������������jkmeikr������yq��teouoknz{xxyz{ukfn}{d]lyxnjlpvwqgm�|�{�{x�y_i{wrnu������������������������������������|seg{�k[glqvooy���y{zoprjeY]mrnkjrukg^_s|~�}x�lYbkdaaekhgrz{{~�����������������������������������zv��sintokjmt|�����������yqffrj``[VRV[Ycvxomnsofff^ZZ\eaelhu���������������������{�����������z{���y{}{t