����OR@����խ��_�VM�\|�v���kjh�>��T=��zۿ�}�<�3Xb��n�����$"��b�t����H]a�Wٌb��q��X'�+Ʋ�2�l���g)|i�8e�bw�p�ɒW�c�b�)�47ͣ�Y���v�76h�;qw�]Gz��5�Q�γ�x����}^ʫ}�\�������sW��w\4�NDs���k
���w��=�r�|�=��S/�j�G�������|�"y	%��EХ�Jh��m�����JӤ��֩kvP���'R˿��$[�������n6��p�r:���S��|`�#���;��ka:-�U�52��D��G�!�y��s�~�c����Ǳ���
d>���t��'cۚk6̄������M�!.�0^�������)}0b�̙³F��mv0��~>�V��AÚO�2�#��Ջ]����uk���~?��Ŷ���+�������tGI���țk��{)�M]4e���#�	S�LN�j�����N�3JZ
�6�l�� �Zxs=>Op�(���q�uع,w��l8Oߟ�J�y��uό%\ 1
/���ա&��ՙ�іﺬ�oM<��6�a�J�ub
�jI���bU�rd�e*���-扲v�k�Z�+�ew��/Y{xͽ�c9�(��:\I��~s���Үm��y�6Ѻ θ`U�.��|sϟ[�U�!�h���V�wG(Ic~�]��%(��N:Er���sq+E��(ݾ\���g)p�BN��k�KIT�}H�oY��7�����;ҿ�>�_�{�@��EL0��{^( ��v��T�P�'4����^�;k9E��0�����������x[���,N�:��ؿ�u*>��&���Ϫ��w��%=����� h���2M��j@F�E��rI�O�>�ø��3��[~�x��L��v&����_֋2-�Unك0RR�ɩљ�b�?Z��I�A��̔ތ��`zA�Y5���M��N
�^s7>:߄�z3:	J:͹��:-x���Y�[��V
�Y�P��ռ�R�S~����;R˶�_	��X���[]�;�g�d�m�j�kW$�'���!J�eNb*�>�V��k���S.����Q�"97ۍt*�}GO�$1��5]*s,4;}3չ�=_�������A���7Z<,R+7�^X��3:���R4S�3��4��;,��76d�����7q�@��7���B���I��>���9�������c4��#E�r�~�Q����������w��V�Z��K&6����p�x��[���q��Tu�WBV�}ˎ#�	\��Cr%jA�t'lk�_�~Ez�F9��#��>�7���Si)������5���1��� \�	�j�*%�>t��tI���i>MBZ�+��I�M��M"b���WI9�|C��޺ݜ�˒P����G��(_��-�e�q���,߇N�}-Τ?s�dQM�@��yu��dq�!��HS��o����u&]�/��n$uh)C�HV���$����u���� �MJ���������q���ԗ����^�?�yˬ���=���W.�j�ܺ�ŵ����Vm����7�O���厸�;�L���%�E_+��u�=��&�$��}�3�8Y��!r��JL��ߑg��4�����!�LvsN������a�{_=�|*��|��;M���@?T���}N��v��.oҒ����]񴲐�W�F�q�P�(]NIY��]K����O���f�F� �}�*��+��A��x)��%�ز+8��ڼI���}}��}� t,��dLYLҦ9��������;+>����ͻ�R�A�����`����Am`�e�k�\-Aw�|v��l?�w*zb-�^󿅁V�@�6|�>�N�1ګ��kצ��Uoh�a�4g�Dty'T������T�n߷��׶����}���я��x�9K�B+��A+�_��j;Ż�7l�m�VH�}P5�Qa%Dqı�TpOqn8&_���S3�t���Շ��������CG���s�ʓ�+7^��U��]��?��vrst2i�P�Q^\�M^\!^A�1�aRA[��>PA�4��[�[My�[��;�ֳjZ�EK�ǵ�-Q����֝�vH��_T��k�ow�����$��-T�OtL�_�&b+����?�H����QV�n+a�wtw~�S���r�{H*�Ri͹�v$|>�_��U9�_�X8"���w�[��X�Miϯ�+��/�I����d�Z�>��:g��B|R��*�%C���w���2��~.V��ޟ���V�~��*�(�I{�7ҋU][��A���U,\Q�h�H�Ty�;[�@�ï^Wi�
�X�P������Kw�)����t���;�>�m�o��P4�≜��؞Hk�R�n���S+���Ȓ���,M�9�N&�Uв
�Xk,_�>� *�-"
n �kI�?!�kJ�������Fp�w4�k���8�1��41x�����
�{M��۱��4��B���>\p�u��5i�կ��%�K�Qtq�<!�G���(��:Qj��F�SF���nq�"�J�/͛�?��Ts�㮾H�c�#TT�+�l�'��_X>����*)b,��,ɺDfwG�k_"���u�nˁ�o��r͛���QҌN�(G�n�>��ᓋ���v�Q!qޗ���_���bt2;�2��ZP���KL��m�-#F�;�%b�Y��q��\#�|�ԕ;�%�@���+w�K 绶�b��.�x�,J�߶5!��n���'�1�-Im��bcԾ��g�.��=�=9�J#LP�6k����r�EN
�z�D҃�����~�ܖ��F#�Sɍ8ƍ `\��$\��s�s\�ƥ]#��{<w������Vt��Ǘ��8�J��S�߻r'���Hy�r�M���d��@Q��P����ۯ��y^��'0:����f�L'��3R��knlkƙ���JH���O��s���D��`$�"���$&0�lA���18��tRm(~�.�=+������]�}��?z����	��RAuzC7���	��׼0���=-�/�)+�����t��#��Hf/�/km�
q:+^���o��ߕ�e�v���9���y��U��y�����ݏ���.�w8�O�jݙ:%0�|�B9�ټ����{ŗ&n�9ks5������H����0��}+��A�ۺ�\c��Z�ط~��-�ƈ+�|��{���҈������~����+$מ�;�j:�p�D*��c|�J�1����G��_4����>�F={���M�#�2�YYx=����r�"�]�ފ�X�(��g�U�[
�A��aPB���8�q �� �p����R�-��!Rɵc���!1Z��E��׃H�ʓ��3 ��QIt�%y��p|�ޣ��w�G�+��Uw!ܟɣ��}`Lئp��Es�e���?�ijle��uS����gd-+��r#��τ�G���idJ�����&{V~V���2�n�?��Xjv������'�{9#���mHbF�'4ZcN:��+S�L�4�:S�@������y%�^����[�z�d��zU��e�M����h�� k\T����(j��y�9��^jϺ��~�J�Q��(�y��]U��c��eߣ���<䅐�@W������Y�E���#��1�e5�t���x�ŗ/�J�d���r�g蚛LG<u��8�[UE(�Mr���g���ݦ�"�Ly�5꘷Z�"���ׯ�%B������s���~�cL��#JoV�v|P�z���y�bq�0*�lC{ ���:>⃷��0	�=v	���:��W���.faK{��_{�;!��`�^�HJr\'�\_'I$�$~��i���l�eXt�:��v��
�0,!��wO'eZ���e�w�e���z�5�w�-)Cr���GQ�"�~��k�k�������� ��"�,�łI���H�ӂ��r����F&f�2��׉��������m�Oo^����h�g���r��^V��c+�<�l#W���:3��i` �ظ�r.��ƙ�S_U�����c�G̿]ߚ+��P�<��Z����?���Nke�%@cՏ����=y���S,�^��^��n�F���l���2��\)����������s+W���;b=v�Yq��g�jZ�;��dj������ړd\E�tی�ł����t���i��d����oeE(?�J�����5�S��Fx9�z���ȋ�o�}�e����f5�+m�D�/��QBE�m�����2��*��YW�~f��n�;>#'��-�/��1ye��7g5]2�bU��J�(ީ5�%�_I�ZNUnkXE��W�Z�ʎa�%�K����Ju�l���d	��^'�����
x�n\�oC,�۞��9cX��7W��G�*��_.[�q@���;��ZU-_��Ѷ�l| g�o�*)u�/S���K�vk����QV�W�����E�j�����㿡n7�mli����V��*��7�L��S��ᬅy0$�+��Mf����]o?�U�t��o�0!�ӷ��ǯ��T��p������-VɨR�ۛ����RP��wO--�h��6I�ne�F�V轂gU�6F�a6׉fF������j���ʼ'V6"��5�&�E��6�S?��j�Rsl>Y9����k> �&�k>JL 6D|�\Z��Mn��v�C���ƚ���f��lGG�ٴayFD͐��M����HC�
�:"�n�A���(��}��I�n����*�1F��c3e�`��*�=sk�e3�y�j�ŒUΤ-j�u����ؓ�i�������3�暃�v��CIa�zW��C�u�p�M���X�� ����\39�S���&*��|��Mh[s���=���`�|�d�rUC%�2瞣�x_}V���u�YHN`K�AX��v�Sa�As&zW3�
����Q��I�� i�q�q���Z�� X�,i�֨�W�{�m�l�m��v���WZ����9��̡�j�s��{��D����!bW6H?ئ��FEQLb�hA��xuVQS�Z��Zq�e[rƆ�ar�F��,�V5䊬-�G��lm�$����T8��D���X�R��D��'��*��M6&���rm�~;0�~=P�qp#8h�ZG߭i�έi߮nW���a�iO'�^eQ��pu�@;ZZ�]�$�tqf`Cv�w�;��VH�