KO;OU?SY�AX_ BYb�E\eDZbD[bF]fKfoUt}`�r����������������������������¸�ā�����ʷ�Ł���9��Ŵ�³�����������������������>e|9Yq8Wt:[z4Uv9`�<g�;f�;]u@`nHfnKiu9Wg6Xd@gn8an:b|:Z~5Ko2Nh6Xn;ay2Xj8br6^n,AX&=H2PVCdm9Yg?coCfu?dy=_�7[y6\v@g�?a�<Y�6Qz8Pn:Vr:]z:^z>d|>`x6Sn9Yw� � � � � � � � � � � � �DBB	EAAGAA956:66;9:@<=C?@DA@GBAGCA�IDC	JEDKFEFBCD@AC?@A=?B<@@>?D@ADBB�D@@F@AE?@A==�@<=A==A>=D?>B><B=<�D?>@<=<89623�423� � � � +6L:K#@Q$BT'H[(K\";H&CL/R]8^n9_m7]i7Yk=]{:Y|9Y}9\?a�?b�?`�;\�:Tt9Vq7[y6Wp9]q;]o6Pf9Zs:]z9]�<e�9]{5Vo6Vd?ao2BF3CI5FM6EL6HN7KQ7IQ5HO�5IO6IP7LQ6JP7JM6HL7IM3EK3EI2CJ4DJ8HN9LS:MT;NU>TZ?S[>RZ;PW�;OW=SY<PV;OS�<OR
;NS7JO7IO8JP;NS?SYAX_@U\AZaF]fF\f�F]dE\eNhr_��r��������������������������������������ϼ�ʸ�ƴ�³����ŵ�ó����������������������������Ŷ�½�ɿ�Ϳ�͹�ǵ�ó������$������������:_r8_x9]7Uy5So6Zn8`t5Zo8at3Yi)CO,GR1T_;`o<^n9\i9Zm=\{:Z~9Y}9[�Ab�?a�?`�;Z�:Sr9Uq6Zv5Vo:^r9[m7Si8[t� � � � � � � � � � � � EA?B@@D@@DA@�645:67?;<A=>CAAFB@FA@HB@GBAJDBJEDGABE?@D>@@<>>:=<8;C?@B@@C??D@@C??A==>:<�?;<@<<@=<B=<A=;A<;A=;B=<?;<<895343121/0/-.� � � � /"=\">X$@T&FV*J\,Nb,N`&ER-P_0Vj2Xn8^n7\m5Wq:X|9X8X�:X�>[�?_�?a�:\�8St5Qm5Uq6Up8Yn8\n8Xn7]w:_~=b�=d�>\v;Vi5Uc=as/?E3CI6EL3DK7FM6GN6HP5HO5IO5GO6JP�7IO 7KM�6IN4FJ2BH�3CI7HO:LR�:MT ;NU�;PW!;QW:PV:NV;QW<PV<QV<PT<PV<NT6JP7KQ9KO;MS?TYAU[@V\AX_CYaDZbD]fG`gJenWt}l������������������������������������ �����	��²�������³�����������������������������������¸�ā���(��°��������������������8Zt7^y9^�:]�6Vt5Xo7]o7]s7_s3Xi+LW2Ud2Wj4Zn;`o7[m6Xt;W}9X8X�:Y�=[�?_�=a�;\�8Rr5Rm4Vr6Up8Zn9[m8Xn7]w� � � � � � � � � � � � B=<?<;@<<B=<632733;77@<<A=>�GBA D?>�C??E@?EAAC?@B@AF@B@<>>:<<8:@>?@=<@<<A==A>=B=<?;;B<=@<<A==EA?A<;@;:?:9<98>::<89:896443110.//-.� � � � $Dd(Gj'A_'C[*I\1Qa1Te�/Tg14\v5Zw2Sj8^j;by:`�9V}:[�8W�6Q~8V�<\�:[�4Rx4Nn1Mi1Qi;^{;^y8^v:b~8_�8`�;`�@f�IgyGcs8Xj?aw0>D2BH4DJ4CJ4DJ5GM5IO6JP6HP5GO6JP7IO7JO9LO8JP9LO5GM4DJ3DK3CI8HN�:LR:LT:NT;OU;OW;QW:OV:NV;QW<PV�?RW?SY>RX9KS:LR9MS;MS?SYAU[@T\BV^AX_D[bF]fKfoXv�f�����������������������������������������������������������������������������������������������'��������³���������������¿������6Vt9[{=a�<^�6Vv4Un5Ym;`q9_q5]o3Ym7^y5[u2Tj:^j=c{<`�9T}:[�9W�8R~:X�<\�9W�4Rx2Mn1Mi3Rm<]|�9]w:`~9`�� � � � � � � � � � � � 
><<=;;>;:A<;644965<88@<=A==FA@GBA�A==�B=<�B@@@>?DBC@<=�=;<@>>?;<?;;@<<�D?>�A==A;<B=<EA?A<;<98;99�;87:899785333110.//-.� � � � L'Da)Gm*Pv+Jm*D^&@N7^m;`u7[u6[p6]v3Yq5Ug<bp<d~:_�6V~8V|7Uw5Sq7Vy8X|4Tr/J]/L]2P`6Wf5Vm;]s?dw<dx;c};`}?`wTtxQs{JjzAfyEey/=E2@F4DH3CI4DJ7GM7HO7IO7KQ6JP7IO7KQ:MR;MQ;NS:NT8JP6HP6HN7GM8JN8JP8KP8JP:NT;OW=QY;PW;OW:PV;PW?TYATYAV[AT[@SZ;OW<PV�;OU>RX?SY?RY@T\CW_DZbH_hRlvf��z���������������	������������������������������������������������¼�ĺ�ķ���������������������������������������������ü�ź��<^t=]{<\�9b�8V|1Jg/KY?gw>d|;_y9^s7^w5Xo5Vg?cq>c�:]�6V~9W{7Uw5Uu�8X|	4Sp/J]0K^3Sc7Xi5Vo<`t?dw;by;e� � � � � � � � � � � � ;99;9:=;;?<;965;87>::@<<?;;C@?FA@A==@>>@<=@=<A==@>>?=>@>?><==;<><=?=>�><=@>>DA@GAAD@@D>>>::@;:D?>?<;=;;;99:76;77:888661//0.//--/-.� � � � (9?c,Nf-Qo.Sv4^�/Pq.H`/KY?iyBl�?e�?c:`z9]w>ax>e|;a8_�7Vy6Sv5Oo2Nh7Yy9Y}6Vv1Ne2Sd5We6\j6Zn:^p<ar:bt;d{;a{?cwTw�Jjx?`u>`vAbw�2BH4DJ3CI6FL7IM7IO�7KQ�7IO
8KP<NR<PR<NT;NS:NT9LS8JP7IO8JN7KQ�8KP:OT;OW=QY<SZ;PW:PV=QY?TYAW[CX]CW]AT[�?S[.>RZ<PV=QY?SY?S[AU[H_fNhpUqyb�z����������������Ǻ�ĵ�������������������������������������������������ľ�Ƽ�Ź�ó�������������������������������������%�����ÿ����ǻ��Dg~@f�>c�Bo�6St1Ia2P`Bl~Bl�?e�>b|:^z9]w>ax>e|<d�:^�8X|7Rw5Om4Rl9Z{9Y}5Vu2Od2Sd5Xe7\k6Xn;_q=bs:bt=c{� � � � � � � � � � � � �;99=;;><<734977;99?;;@>>�D?>�@>>�A==�@>> ?=>�?;=�?;<><=?=>@>>�C??A==?==?;;?<;A<;>;:=;;<88�;779771//�0..� � � � A">P&@N3Vm1Yu3\{:j�2Tn.G^8SdCl}Do�Bk�@e�>b�>d�Ai�;a:`~9_}7Xw5Su4Nn1Og7Xw:]~:\|5To5Vk5Zk6^n:_r;`s;as:bt:`v;a{=d}Ks�@f~6Yt6Xn;]u4HN5GM5HM5IO6GN6HP7IQ9MS7KQ6JP7KQ8KP:NR<NR<OR:LR:MR:NT:LR7KQ8JP:NT:MT:NV�;OW=QY<SZ;PW;OW;PW?TYAW[�AU[@TZ?TY@T\>TZ>RX?S[@V\BV^AX_NhpZx�g��x����������������û�õ���������������
���������������������������������������������������������������������������(�����������ü�û�ö��Gj�Ah�@j�Hv�8Un2K`9WiDm~Do�Bj�@f�>b�?d�@j�;a:`~9^}7Zw6Qv3Pm2Pj7Yy:]~:[z5To5Wk5[k6^p:`t;`s;as:`t;^u:`z� � � � � � � � � � � � :88<98=;;>::512623866=;;B@@A==A<;?==A==D>>A==@<<A==@>>?==�@<=?;<?==@>>A>=A==A;<>:;=;;?<;?==<98;:9�<98=87<76;77;991//�1/0� � � � %CS*J^(I^0Sj1Us4[�8e�5[u1Ne1O[FhtHm|@izChwBj�?k�<bz5Vo7Zw;^6Yv�7Yy6Xt5So;]s>dv4Ul1Pe1Sg8]r?e{?i=g}=f{:^z;`}?h�Cl�Cn�?h�<\x7Ws7LQ9MS�7KQ7IQ7IO7JQ�9LS�7KQ8KP:MR<PR:MR9KO:NR;NS<NT:MR;NS<OT<OV�=QY;PW<SZ=S[<QZ;OW=SY@T\AW[�AV[@SXAU[CW]@V\@TZBV^AY_BZ`CY_Spyd��~����������������»�¶¿�������������������������������������������������¸������������������������������������*�����������������»�¶�����=`w=b�?f�Bn�:Zv2Qf5TaIlyFl|AiyChwBk�>h�;ay4Un7Yy:]~6Xt9Z{7Yy6Xt5So<`t=bs3Qi1Qe2Th9^s>e|?h=g}=d{:^z<c~� � � � � � � � � � � � :66:76�;87423533866;87�?<;@;:?<;@=<A<;?;;>:;?;<?=>@<<>:;=;<><<@;:�>;:><<@<<?;;<88=87?:9=<;;87;97;87;77:76965�9771/00.//-.0..� � � � !CQ(J\,Rf-Sk2Zt4Zx6`�Am�=e�9[u4Ud?amBfrAhuFm|@j�<e�;_{5Xq9Yu;]y6]v�;`}6Yv6Xn8]n7]o2Rh0Pb5Wg?dw?i>h�<f~=ey:_t;ay?i�@fzDm�Eo�@h�;ay�;NS:MR9MS�7IO
7JQ9LS9MU7JQ7KQ8JP:NR<NR<PR<NR>OT�ATW?TY@SX?TY>RX<QV<OV<PV<SZ>R\=S[=SY>RZ?S[BUZCX]BVZBUZDZ^E[_�DZ`)EX_H`fNgpRmvd��y������������������������ÿ�����������µ����������������������������������������������������º���������������������+�������������������������ÿ���<d~;d�?i�Hu�Bh�;\u6Wf?_m@epCjuFm|@h�=e�:^z4Wp9Yu:]z6]v<a~:_|6Yt6Xl7_o6\p2Ph0N`6Xj?dw?i>h�<f|=ey:_t=d{� � � � � � � � � � � �  955�965:66401511743<76?:9�=;;@<:@;:>::<88=;<><<?;<�;99=;;>;:<98�=;;A;;@;:�=87;87:76�:98:88977�8661///-..,-/-.� � � � �'M_(O^,Uf0Zl0\p8f~7c7a?m�<d~:]t8Zn9Zi:]j?coGn}Ag�;_}8Wr8Zr:Zv;\{6\v;b}>e�;_y6[n�5Zm6Wp2Xn8Zn?du@l~?j�<g~<ex=ew=d{?i�?dyAiyDl~Cn�;by?RW>PT;NS:MR�7IO7KQ:LT:MT:LT9KS8IP:LR=OQ>PR?RSAUWBWXEX[�CX]BUZ@TZ>QX�<PV>RZ>SZ�>RZ>QX?RYAUYEW[EX[EY]FZ^F\`�F[`FZ`QgmYv}c��w����������������������¾�þ�¾�����Ľ�¼�º���������������������������������������¾�þ�¿������ü�·����������������������������������ÿ�þ�¾>m�=g�=f�Cq�?h;^u:\p8Yj:]j?eqJp�@f�;^{6Xt8Zr<\x:]z6\v�<c~:]v6[l5Zm4Yn6Up3Vm8\n?dw@l�?j�<f|<dx<dt=f}� � � � � � � � � � � � 965955�9772./511955=87<98�;99;:9>;:?:9=87:88;9:;99<98:67;77?:9@;:�>::>:;?;;>::<88?:9=87:76987:76987977743�644645/.-�.,, 0-,� � � � 3(M`*Rd*Tb0[f3cq3fw1^q?r�>l�8`|8f|3Zi6Xf=`w5Wm1Ui6ZlGk}Ce}:Zr2Kd9Zm=_{;_�6Wx:_|?fAj7[o4Vl5Wo<`�