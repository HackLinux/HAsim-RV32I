���2�7�c��+��܏������%
ǒ�%oW��8U{����Kc�(�-ˀ�q�,-.k{Lpo�I3�y�F@�����9��м�L����.(�"bt�02���+1ʳŹLZwyƴ`I��l��h'Ra�>�4�Y������/;�j�
���V���y�Ur�K��r�=�'��m�1|��\h⤡��hS��"~u�r��*H�0�|E�3�UT��@T�G���\��TQ-�),t�x!�Q�-ܺ�:E,�F�#���nvPd�������t�t{ӄ~]�o3>�ز���2t��0QnFSPÉ_5�+��c$̯cX����9�'���tP�&Z��ςXwނ�!�Ǚ}b���߻Ҋ��������3��m�H��g�c;<=�3XfgŞ�^o��.�+�޲� ����8r�Ho��e��A���
;����p�U�/��4ܨ8܅�jPA�4�B�;�@M=��vi�:Ga�,U��2�:*��C��B�P��¸I��l?� �Ao/��5��]g^�G*�eFW�dE��}G���K&GY�.�.`?���L��s_�boTv]�i~;�B˥��Ƥ���̇ag��m�qWA�Z~�Y��t�~5[s��N!pN�?���/�0.�Î��qo>�(�Ry�i9�J��jѼ����~�J-�����ޭ����7�wА��F��Ӛbʒr���*o��G����@��Z�2��orA2�Д� �m�sG�U�e�1j�����p��lpZ��G�+9�;�g�;`����� �N�����C��A��ͯ؄����a���ݘz���5Sq�)Ɓ�66E9��W��[[tp7G�Ej�n7���2W�Y��V i�����y�Έ0��&
�.�6���s�/Y�h0l��SÖ�,�A����yA�`�F��_�F[nd�mDOV���t��Cq���@p�9�V���F�7r�Pm�e�;D����4g;1W]���gX
(�V�/4&[�@Կg> Ó]�n�X2��2Fv R�m����>tK�eî��-@�cZ���${
o���D�)v�,�K
C���
s�#3�UE����zn`��n~���U�R�R�
�-ec��fn�-�k��k��q��+#�U��d �"&�䪓E2���W%	�eW���7ZHCXOBo/�|��|���a��95��� �pV��e|T:�T9������}[u;g��>�l��ƹ���q?U߀ j @����8((��g�<���n3�I�&v���;a,("ܦ��hNU�s((�h�r!GQ{��j&��:���n>�`���'�d�!b�����͑�e��;0�=�^�K�b������%^�������:~��ʥ��H���@���p�t��0k� ���R'"#��e�V��q�2k&�Rn��_�EdFؠ<�y1��g�*fi۾���GuǜR�a�k�#7��l(�~��, ȣ����Ƣ��i�6Ja̎ST9 '��D5�f,�@ѣځŅ��|$������e�����}/@%�j��<���i�u�R���E�|�HN6xV��P>j����G �o6���!�s�$7u�5��f�"��u���2ùwsU�E�� Zɯr�=m�=����?��T�}֪��I'�C�o�1�k2��ϰ.!ύ!m�*6�b6gA�X��t�E�c#|_x,5ê̞k�n0cz����-r�M�Ğ�~$�ϕ���`��My�����|]�w��k4���w�h�?�ɪ��@��e�zC���D^��ߎT#[���$"��xD����^?�O>�h=4�.����V�I��Y��.E�g���m&8ϸ�EG��<��!�R[-F�J	�>�!��K���56%���n}7/�I��al���[$�����-G�߫_#^U�,�\����%�ے��f,�1�����-�{���H��=*��ѧ�v���Gr�j��(��sÕ�)���!&������<�%�7�����]�%1ͤ0c����v�r.@����w٭�T[�Q��&p�6���Ɩp�/�C�@`�����{��S-��9�&�b΄�P���rٕ:��<�R�+���C?#o�����'���7��9�rރK�����"԰����r����o1%> ���nkn
T��C!�y�ZZ�Ij�o���nb_�q���TTj-jB"�h�t���?K��u����ғ�*��BB�bX��p��������/������)��y�+7�*�T���n@2�Ģ����ѧ����m;)�3�	�7n$�j?+":�W�0s)�6��A�4���e�afa�ŵ�B��PFR�e�6|���Uܫ�6�>̔7�XF�i�+,�KP����&h
�/��%�V�F�q;��PA+#�� �s���fi�*~a�YŽ^�mkL��?�f�#�I&+