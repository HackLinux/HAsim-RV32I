oo�oum]mu����_N CG)G)DG)7G7G77C7CCC)D)GC7D���b��c�������            ���nª����ttttt������������������0>������0�$$$$�$A$�$$���$$$$$�$$$$,U$�#*���^����00�r�ь����x������UU�U�U�RU��tt����c�oc�W�oo�o�o�om�mui���_X C)DD))GGGG77777CCCDSGD?CG)C�[�{b|���            ���c�����|�ttt��R�  ɵ������������}����0>�������0$#$$"3="<"=#######A$$##=###$$*��������5.���w������p��ȯRU�U�URR�UU�tt�g|�cnuc�Wԋo���o��u�]m�����f� )GG)DD)DGGG7GC7CCDD)D8:C)7��_j{���        �͞�ք����Ԭ���X�       ����������}}ƕ���52�������.�&#(��������50���w�p٢����p�UU��U��URR��tt����cn�c�Wԏ�oo�o�ummmuW����[� ��DDGG)GG777CC;CI))G8??GD8s�q�{b�c�   �͞ۄ����ѐ��������            ~�����������}�}����0.�Ծ���('"@+,,,,B,B,B,,,,,,,,,B,,,+,++,,,B,,,,,++,+,+++,,�#%3������00ɍ�������q�e����U��UL�UUR䳵t��|��luc�W`�o��o�uummu`����_� D-�F�DGG7G7CCCCDGGG??8:��Ncf���ۀ����uu���\W������           ��ě�������������}�}ƕ���0$�����(B#                                                      95������0#0����v��������H+U�UU�U�RU��tt��|qͅ��xWԏ���h��ummu`����p� D�-��-�)7CCC8C)GGG?8?2�����c[a�b�n�������}����           ��ϫ������������������������|���.0���#0%8                                                      4#5��ز0.0ɍ���v���p������JUU�URUR�J��t��|y�k�cͬ���hh�����uu��z��p� C)I��IDDD�8?CGGGG8?