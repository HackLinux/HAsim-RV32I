��:�Y	~wz6>X<U���4����O%�Þ2�����]�v�ɫO���U���s��?0�x�k���<�a�t������7N}��;�j0m8܀<�!j,��S7�5�w'�&��C��Y�Xľ=;�6�(��~�q^�>��빵o� /���
u��Uڐ�n��%�m_�����Dg�.�D����q�z��9��ݴE+�f��d�����=��:v�N�8�t���G��ğ�C��O=��R�0�C}����~��X�j�,�篌�����I�_�g���{�:�e�0�?�x=?����UaPP���8F��\�����³яJO���_�i���f����F�:)-[��u� b4{ăs}�G�f��0󘔋��\}F��{�ݣ���q#�'�i�DTR=�5�z(y`k�Hq�L�S�������Z��&xҿ4u�,���X��@U�j�v��Y��}�Mʞ���oNf��b�6�%�Լ/��}�w�fà��%�T���_�'LzG]�n��B*k�lA�^u,���D[�+M���5����~l:��dFa��e�FߚO����dz��������S�߳A�:| 7$�j�S#)ǂ�^~L땧��`q��<T\6zmH�S{@�6R����K�Ʒ�ͷ�hWuW�y��v8��lH_�Ùޡ��|�p�	^�5��8��E[i6�hu��`������[��#����v����k+�^]/��U �kG ���f��|ٗt����cӥM_�������L�	�.�W�:����i[�3V�As��'��G�|�3k>Jk�ܦ�Gl"Ԭ�_^U�0)����?0����UY[�V�����ċ�/i|;���\5x�z��d�$[�EO��ԗpj��e���F�wP��d�󻫵׷q��}��U9��4*�=݆N�
~_�x�����+R�g�D������ωpE�8!�ڇ�\�ܻgS�鶗�+���+ox�$�o�d�S�;��eP�CAo�
�O?_�+�;�p����f����AǶ}+Ť>ݶ��fTS����fr� W�|���&��"<�m�G�fѐɺ�1	��:����"���H�;p�f&R�M\�ۑ�`V�:��ᕬ`�{��1Z�yBJJ�ѫQ����4��᪀�_�k��[\��z8����`�7���Y��q�G��擉�>ޫ�Gm����æ射cF!iP�S�E�ٽ�b��H�g�q]����q[�?z��������fJ�7�i�C�-���+��ڞ� =Wd.����1��;Y�: f��z�ע}�1�ъXc�����G/�#d���<o��.����?�m1W�]��ģ%#f�k��_K��E�~������^�}���:�ޞ��`g7K��K���y���e�~-#�>�w+��q��ݝ�ͩSKf:5��u?�ſ�a����H����]�~+AOq���Re٣�J�������k�I�qO���byġ�'�ԁ)�����n�&s�B�t�%$�m�lE���h��4׻��䅉�J�z����	�NkxU5ؿ/޷� ye���5Jj��;@��"���kB@Ȩ�j��Jۨ1-QL���>��E�C5���ݟ��$�r����t��u:1u.�a�wtx�UVlA_�8�Et�n݉�k��MC桨�YJ?��P����CE�j�^Y�@����}�]f�;k�0�4Wo��amnu��u�R��͡�U?~���LY?C���!����}����J�����!M�I�E:�\�H�ل��i����=�.�sd�>�Ⲭ���3W�й��7�v/�O��4y�훼Ey�x�Ef���fޣ�g�{��-��>x�:3�V���� 9�j��YBʨ�����W=���n�*L;�>��k�8�<{��R���x���,��.��c�u��Ð��L�=�O�����j�����#���~[$1�ͬ=�u?�\^��e<b���+��e�ee�1�9�%�oQʋ[��ղ�q`�o�M����t?�PY�����8��co8��v;2���u�tu�������Uկ�)+��{m�W�q.�t�oZ�Д������>���ȞC�=��:���ec��Q��J ��ĝ>)/r�]1Q4`��Z���eq� +ַW��E��Yڷ�dJ��y���,�uE�]G�|֖���=�ۼ���5���+�x�~���3��g�|]��H_���5_Cw?nشh�=�`�D�W�]�I��L��̲^�4�.�>%eRn?�&|���݈\��֧5�u<λ1��{�D�K���潵�L]cC�,���3�U�<�)�nH��u�SJ�ͫۢ7���5L��IE�򻾘mzf��S�Ώ�R�����%�r��M�Xi�;5�l����p��E��U��9�ZĘ�u /52�ޓ���i���f�G��͈£b<U3&�x�/iβ����<�aÞ�
һm���j*l��KC}���Iם��k~^#�違��|7�N�qm����<u]�.N�[^�����`�M���dK>��\=hѼ��CQli�E�L�&6�d?
h��9���R�K����M}����G`cn�\wB�[���W�f>ۄ�x>�ru���y�dՇ�M�� oh���_~�~c��U@�V�D���K�zF���|��!�.2����f�I�z�g�fQg����+�����'M���ĲNF/n|q߯��o'e��T��՟��Z����!�k����C��OVm�[�h��AC���L�6��|�)�c�Z����>�f��w\r�au�����B�����.:x��j2Z^�}��U{�~�	��Mu��rCɁ�aب�-
���g5�d[�'Js���ʝ��c��:"�7��˟O?�{���D�C�w+
�������Բ��7��^׳3�G��y���U?���_mW�,x��<�h������"��^Z�����ϑm�j��ݧƖ�L�3�X���V~��bO���!U��6^��9����βk�W̿ߐZ�xy�U��ay�Vx�@m++e�f�0���������J�I�Rә�)_sCo�ܚ$<Ys��2�!��N�7���:��&},�S9��&?t{�w0�{�"�s��d�x�n�>?�c�ኟg����߲/W!����=]y?H�����:�������]�j�?�ڸ���56w����2�ջ
8r-�e�������frP�^mv]G�ls= t�M�A�/�}w+Y�0�[3���ܚ�.ݭ��+�mu\_���R�T�u�}���͵��z.5���\}/��I�*�������M��4���q�Y�I4��G�"����OXp0&�I��Ȯ,�U=�\�4��[���<3���o~~�x�Dg���6��}���=\~�0e�Ӆ�Mnz/\4���~-{E��஖������~n7j�����_����{~G�X��������'nu�y6p��>�J칥�z0^��F�c��u��&ml�3�N�}�@֨���V�������Y�By����r��R�8�ҟ�T�nwax��Am%��1��:�+�x =0���yJ���PB����j#گ��v��3���m�O������.ސ/��#~\�R~�}��u�c�����;H�7��f&�l�n�����>*� &յ�x��ǧkmx5#S��\A�$��^V�x�&��C�>��������.RGfOqT�#���=�U�&ÑV<����餒s5��f�}�춗/ԫ���k�rHG�n~V�d�8�����qD=����gv�z	�)�rM�b�^�����*�c�G�궠�n�Y�R��l��k�#k({&�������b
����=opָn5��L.��^��@�0њ�r4I/��qڹQqȸ����W�~�}NB�� ������%����W�e�oXsv4L����� �(�!�7���3�t�E�=��m�#����W�4���z~p����	|6rbu���2.��nw��B���M��oS]�\�;�������J��[����PN��~�M+'��ʨ�]7�fV���gn��X3���̣��&�F_�������Q���Y���G�|�5"�_%^�v���*����۴�?U>����WA��"�]�ؼ=��>�j�i�<�Lv) �Xն��=)Vy�SsF<H��*o�bO5�ؖ�_��f�TӿQ�{/��q�����~�sZAH�{ē�ۃ�ΰ��y�k�f��3��������v�s�97�g�^V����]~4�$1���doיt�}�V)h-��m�KP�)��.߬�3��#U�5ǍR�Gf��Ǜ�Q�CQ>���y��q`9^|�l5���d|'�Zu$r���I�� �����ʟ�3k��?jk+U��c���b�免~��U��U�[�}t�Z��#aV�����p{s��HuZ�i������/0L��d�#�WcE�7�}k�y��Grׄ�����#��%�O<Q��%p7�r���\[p����q=#�l6���<�^{��3�����gdM�̈́�b�\�Zmg�Tk}�V�#��+`�<�G�M�	��o�I?w����5���]��>/�܅4��m��g�규nt��)����j��P:Y��H���(M�SC��/L���L=i��}�T��^�)]�v.Il����C�0LYUU3�ݮ��'|ۧ���AG�T��0��}�jC=Ivt]��'�G������֘Pkc�T9�F�k�$s���Þ���n�͜yN��8�z�W�F�"��������Ǵd���3��lg-����Ճ����2��B{�N��?��h�K�C!}�x�ħ�x�5��f�u\D�9]b�8��^��^ָ׷yi'7�������r.�XE���u���=�Ҧ���l{��J�[�}ˎZ�q���_$���l��YX��󛳊w�F��lܰ9�u]oi��|ԉ�X�m^&aKK��C7^�4�Ӿ�7{��C��!^z��d��i�:O��z��C��w��:���O
m�=߂>�oy�dO��lW���0���c�3c+��]���h#����^��
uܾ	��7v�e�*��]:g��:(����ײ��"B�3"Og���a��$O�K���n/����,�����Z�;�|(�y�=�"/Hh��TqzYI����HX8�;�z��Y�czmG��p��)�ʀ���Hz�>x�>�{;(�R�'!���Ⱥ4㨔����g��:5v�qn��`O������C��1������*:��V1�]�K��Po7G��"y(1���y�z��"����59�_'�o���f�׆��^i�e�.�ݸ ZO�Y7�����!��/�و�'޵M����{WuU�_n#`���[�D>_�1�V^��ސ�$3	v��|�o �ua}�r��TB���{"�ѯu:�K��.����0��hk/�RhI�xD-q�c�軵���Ʒ�W��~���u���)�{�ݛ���Kӭj�������,�໑�VIU��u}�ɫ~�Ɲ���;/�$��
�_
5|���[��*����G߀l�����\.?3�!�#����&��:Sz���������1�T$�B�+uot���J� �~���x�mC}���l�ty��Qܴ�7������Etŵܼ+�����������Y.�W�[�[b�2_U��y�C�7�~��E��؜=������,髺�l���x�2��n���	"ו�ކ7�F��׹)�������Ý%�m�%;��[fF�3���e�w��m�V��dE����[�w�Ku����!w��_
a�=w*K�?я�թ�g_��Zҗ�dU��{PN4е,�[�,k<k��[�%�A�=�.?
�ej9���39��b�nL�������u%��s�MU�'��WZ!�ۘ��M��zj�Q&��8A�0�bhm����_�W�K/�7��tޱ��g��,1�֐]9o�|B18&}�,o�I�7�FS7��a���X����[���]��q�z�^q�ԇ��_�i��M�dg���p�Ҽ+�k�����7������usCǅwڃ�k+�B�q׎h"wȓ�����;*Yڸs�Kmk	�y1���/T첗�s��>�4ۻ��Ӛ�l�zq�F�i �HIe##:��;!���=>WR������jN����G��i��;��ݱ��{��k��'�Zw���
����Jt�\��--hn��橱	�����岑�d�L��Z�f�C�����Q]Aw`	EN�5i�˿W��m�}��DS��2gC�]6�H+D�y3��%ᗊ�g(,�w�o��I>Y��xw�p�Cz���6i>{�ҧ���2�/�򚃅^[��=�Ml�#��ъm�;.,�1�6�nK<c.<�����f���g�څ�v'��/�Z�W�;���m���p�{�Ǉ�kO^�S��2�)�K�	�X�.r������x������c���I��ZߞN=�η���&W�Jטn�%��!��QoB^�\�K�^P).jg�1�%kZ�|F�~���W���oK�k6��ͥ��F����6p��Zdv4���AVb��%�Ǳ_MaEzЇ'JZ����F��O;љ�g��/.ˀ+I��]e���,^r�-��w�l�����>���:6D��p��{��:g�dƬ��(Ի���I:����(����uP�/jK�|2�W��j�,y� J����`�Cobb��wD����4�l����������qW�a���ֶ/�����j��b�7�\a�9X�ߏ]��_$N�ju�fo��酧߼�>T��NڶVז����}����/��F�����CM�{�n�����y	�m�L�W�G�c��'��� �I��[y��:U�����A�����:�Ǹ����<bjg:���dw��Z�[�����ћכ>U��̕Y>�:_t*�@��)g���X����]{g�t/2�͠�M�	؆�[qy[���t�ÿ\q`�c��&^�{���w �ҺCf�����ֆu�;Fb-T^��M.�꿡���C��GsWt�#���{��Θ4�[C���	�s�X�*��s����Gw�;΢Q��?����FsX�I�������4Cƞ#||����5ko!f||�u�b{g�~Ӷшa���:������W��Gw)�&����r]��?�`�?֊�m}�t:����v�7�k^2���S�u������v�&�O^���~��%�w,��ej�I�~�O��w�RNm�lq�>��B0�f��M���֞wA���9���:r= ky�buAJ���=5t혒�N�E����N�_���p�E�p3�*������v��+u1{<�rJ�xg���^#�2����9�ڽl�2{��zj��͜�N�}����������I3�ڮr����q�Ǯ7�|0W��J�@�L:��`��â��?���|��^>�F-)">�G�^E�;1��;>�ekʬ���q����+�3s)�-/�L�lwd4�`�C�l� ���KF�l���^�_MW��8B^�Ej�k���]~���Ğ�3��8������C���Ɋ�z�}~C�(�G���i&�,3�����������|�;������`�c�;��3h͒��yU��˓/��vD���q�`<� 
vc!xp�n��_��>.7U��1���}oL���V��3�M�3q5.FR�\��O�!�Ȣ�[��殂�xܳУL��U����i|�7�s�����3mq�o�B�7w�##K�d���g��LN#_]�r�l+����#��\4�߆vU����N�P����ֆ�v������W�>��v��e�5�Z�jJ�.�j��x]Cb�/�۷�{�EOl�p����)}c��ܔ�wq����b�����x��'�0��
B��q����s����_�Ǯݾ�`�$2��[,\BL�Z@4b�����6:>y�}�{���|�Ǉ�&u-+���n.;��r�9��xyu�����y�n�7R+��������Ǹ�w2m}��[+wݬ��_�N����m0&_#<�76��M'�n+���Ng�4^yY�h ���;��jt��^z�h�TEf�����g<��~�͘3W�x�T��)WjЖ�j�Fg���S�x��6����۳��#�R��W�䜰���߼-�wv�g�_�GyU'�rz��H���x�R���a'����Z.��s��Q�ݦK?��־]�v��a#]� ���^v4њI�U���  	/���X���Q�Ow���/� ��5��S�AN;KxFa����+/�;�Hxo;��|�}ܽ_�j�w�o�G��7=��)pd�8#<��S{g���0�,������'����A��;�W�DZ@`�>��
���>��s�)���]����O�!=��H��|��z�E5
���xS5H���˦�]�Sv��C�s��%�h\Q���"�ؕ��{�l�+a�V��(�yI��g�"��r/o��|NI�J2;�ǈv��v��:�v��W�5��q���]����9f���9Gc{����g��6��H�,;ߒB:��a�.�zi"�̍2R%�İ���F]��D����_Α��7�|<!�X�Z�~5�3u�X���
}t��1R����,>��Q� ���Η�	3Ϫ�����+��S�c"��#���U�/2Ի�D��g����rg�q{�?�����H�;y���sZ�^��_�n�\y}ܳ��f�ˁ�Գs*�E@+zy�]��T%�|[˄��(2�K�i �~�����'�^�&BF��}	:�1k$t�e�C����O��×gD�0��l�h�)�a��Qႈ��U�1Ŕ�O�E��A���7�fR�*�\�Jy~�'n?�}�`���jTĕO]���_'��t���=�*�9&�x ����z
p!3jC\C��B�*}�Pt�nMC�b5~�k� ���%��oM'��u����@ ��|=��r�s�����U����`;7N�w֔M�� �AW�E�:I�;V÷Twn��E�^���s"떕�\�zŁ��}OC2M����ц������Vy>��g2uK�=o��(�	:���KG��mK�{<�;�e��Vc��j��s���qi������Bªt-Ŕ���l��������7hǞ/�4�[EK|�#����rڭֺڦ�NR�=�z���Z���gc���{�ۣ���"4�(�����ˋ��eRB����گV~X���@��qS]K�.��ҷ��9�$�㾫}�Z�_��ۢ-TgGbQU4gvO-�[TM���1�F�/�*�Ⱥ0�d~E-����T!�&���>ݷ��~�{�������}���{E���v����or���I����uU�ww��#G�=�,�-���8T����o�&_^����P��!o�"f�����o����Op¯(˕�0S������\���s�A��'��E�~���e��c:��+����]��q����#��oeϟLR	��P����k��/]��a��[Y�'s���>���=���>'�S�s���s>��ͷ��9�����[#K����î㛕*���Ϥ\���0�Q;dQ>�=�ȬN��ٜ�yv��)�����K����O�AS�7��`�a2��_�Y�Ɩ��in��=x��0�\+��5uul���oEG[C��%	i/_]zU���7>���������a)�8��y��R�cWF��!�U��:�?�^�a\��{�G~�y�d[Ɍٗ%70?Ry��;����N]^�6k�r�����o!�u��8���꓅�����
v�`c��9�!0#b��M�������+�`=��2�'3�wnp~��q�<5q�2�|3�f��q��P��N/�
L�s���7:�
�f���E�lJ��[�O]ф/+{�B�.ٽ�C�����s3SW�����&nb���c&����ǚ����u`=q;C9�mQ�\���\Y{,$�nSl�ٗa�ǎ��*S5N_Ut!��zch{г����_��c����W^�	���>�!���C���Ԓ��w{җ�WE�G�.OO�=2%��GU�N4^��EQ�1y����wڶ^����^����<��;�`ݥ��I��cEԛN}�}�IR-ֳ����Kܺ;gvf^s���X�\[�~M�Z�xPA޼V�5s��S_�{��\h�އ׃�������v6Q���~�|�q@]k�Vϗ��=Qro�rnI���&[/N7:mD}��t�����y���P֗�I�\�/oܲ��r�V$hΪCzV}6�8)M�������~T�����&G�	B��+��>rVp�g��6
�W�kȗ�����J��\|��U�dS���?_�����_1m^;.��^�=��7�8 ��;�����T�;�@>�:}&�?��tĻRg��"�^9��˗�?{�ح�y�Df��e�Ve��[����6?܏{ѳ�֤�F�~�S�U{�\.f���n[�i�����KbAÈ�J�[�)�	u_��a��C�^9ߊ��aT����S�V�9�c�����R��[�Ae��[��c�F��������YS��5>q/�X�K���O�}q$�ð������dq�S���E������>es����s4��+ω������ҽ�M"�8t:u�����T(�rxTf~��zlˤɳp�KEI����ꗗ��������9t.1�t��:RĄ��q�է��O_��w]�X+�{��޸�Y�����|�E���7���s��A!L��N�J�va�a^g�I�
����d��g�N$O*S}Y�Ysa���M�p���ת�,��]q<����o.�iK-ZV��o�Iʷ��~[,�_Y��?~5bS����C�զ��'�D�++�Aw������w�Ϣ4�Bz���opuM�=�7����U�εO7�*�]Jz���z\0�19n�		1{,;}�YcN;X|Z����]�~�b��|��}Jc���]��m~Y������#��ȓJ�}ulC��:J�r�Y�7��R�Yu��C[?<˞ث�t�x�������[l�5���o��^�+��߳2��o>�x����݌G�S������˧�;}!�������]�j!���]Ѻ;�߫7��;:p�y�z2��z���p�"]*���&5�H<�8?��;?rt}Y�~̣�çv�-��wJ�2�&Syv�Q�r�,���QCM��G��g.��yi5�D|]Q��8a�o�dC��Ţ0���q{�����|5q�p���K$إ{��}�A�	�W}�ڤ�c�TS��j�Ӛ�Y��)R<5,�P̇+s�&�]�M*u�wj��5>���ڃ#�� hW���s��N��lhk\RÆ�����n�%%�*?]�;�=%����:�P�y�4kuzյu�*�.��=�'!��vM�ؐ�E�w��|t�|�?b��+���_Ņ�A'�*�n�y{p﷮�൹��e+�4,�O��Lu�d9��=��\j_�o$��'�(ߒ�"?�v�㧁��ް����:�җ��Zq6���Ӈ�<�����.X'L� �$׍�ro����nׯ�1&�2���:�2�7���SUK���&���zO�D����vnL�r~��j����'�~�Iv=���U���]/>����b� �ΆU�L~�W�0������/6�QI�ۧ���bn4�o�#u���ٲB��2�Ș��~��m]%,;�x�6���o�\���fե���7�£Z��������;6�Ћ�wW����`es~'t����?����e�|�ы��q��WK��뿰WI�?�6_l�s5$��2�^|�Nq�vWSA��:�$��:��Ѷ����+��.|\4��w��
�4?�������\}r�~���QP{���7@������F�F�9/�N����=�+6N]��C�c�Cb�_��D�FvV��e��R\N�~�Q}�{s��-����.֕�~����=��y�¯d���{w=��~������3A����=+����}�A��Y:玆9<�:�:?�i�W�̽�S
���x��c�2�l��v˽�+�;��2��C�*}���a�c�
�1p;l%�i}��Î�a����?�an�j>�gh?�[�����(�8������:.̄ݵK	��ZC�,p��t���7ۆ�Zx>z6������1���[������md�|�Ȳ�����~��~��Y-Xbd�Β�n�T?�Q��Ή�3>�Z���nͨ���%��T����u�+��w֮xs5�ԅ���rj�d	U��#,LۋX��t-w�XC�P��y<�k�JY���k��i2���Ұ�����n{���t�ﷇn��kn��HT���n�w��ր6���;��=��-����}*�=�)�R�����y8v"o��F���M��Ҡ���S%�җ��KwgO<����qu̾�'jZ��/�Nes��� ;;�}S�7)��r'~*`kHf�����lh"p��͇��`�Ǥ��9&N�b�d��d���_���9Y>��qc�5>W������:Y��&?yܒ�[p$)=�trb�c�7a�ovGu��Cw{c��铢�鼧6i�\s�gwtL.�U{����!�Ï�2'��ҘJ�K�Ҹ'��YЏ%!Se�\��W�n���ѭ���X�jlbff�������UK�I�-�|��/M�l_#ʕgz;ށ���M�m;�^�mG]1��R��v�;՛��|/e�0�p��ʟ�	2'��c[�J.�/�0 +'+!Aץ�0!�6F�,�<q cRj�I�Ҷ��ҦM�c��-��u9}��6����mt:\��#��N�Ը�ȯ��_�қ����I.���zL���������i��^�(`���k0��Q��U~�x��Mwu��9������:�7+���~/9��t2	!_2�j!)�TϾV������u{	)�փK_��
�gfc�rВ��Br����A��!Q����ei�y;������=���lw�f�D�c\�c����+��=QW}cH��y�㉟W޾y}��1l��Rծ���s�;�*B��x��7]��y�ea���]u9.����,��"���G���j~A1�/�(s�u�nj��Dd����;�֦ڪ���b���5�zQ�c���Y��k��xf�ͱ���?���pu��ԳuӢ�g�+;�
�߯�|S}�`r�1��obB�o^���������P���s�"Q��,��x��?7���s�&�^ә�g��;��6&��b��&�gq�#:<���d,�8�.��A�L�ن�UO�O�P�#)�"y��^�������OsL�~DV-O��o�<{�<���FԯTc�E?O_f߰�G�7cw/��v2X���?3�U��~1�B��q���sر�拄<�O�N�� a@eD2X:��ؒV�/�vk[��mC�5��ͼG��'��v]O���,C�)r�(@O$������莛*m�7Xtլ����F��e�S��������ߘǧ���\�:�>9�Le�>���0�i;���g{䷖N��ȟ��&x'#;�?Ĉ����:X�{��p�ao�����gS�'N}�&.m�i���i����7�����xX�F2me�#��2��V/K��\�y���������.F�'�u��>Z��ry�o+�R�F:�w~j����Ԑd�_?�/��>���Y��l���C�}h�s���&�HGS�g���4��aV-o[R�훎?ۇ�.����~mSo�wk�V���I߫�����!+�׹]����q����o���s�O�v�&��m����_�U[��;��Oc�����r����m+�Q1�C�OkG�M��J;7��dՁ�6�S�<�uU�U�`��?�ֲ���o�����+'v��.�+��E��d:̛{�+*8Q���&��|���������g���!\��?5_��"�t�b��03��ev~~������Κ�u��?kP��)�0b��c��Φ��sᲬ͠*_7�����t#��2ˣ{�27�W�7ߙ`NK�ro_���8�����L�&yu�L2D9�q�;�7lv�Ġ�ƺ�_Z�����l���G����"��^$����!(�7�k��� ��i�N؋�Զ�D����h������P}ns���s7�|����nzj�����	�cӏ�������˧W�YS����	3H9H_��a�\g���Ï���<�������S�v��7���eu_�p\��4f����;���wey ��q��U������_��z����U�}Q����5� [)?o������;&�}��L���/�q.�,��\���n­~[�>���޴�<q��g���{��G�zI-�*�!���cz��<��>5��~�����Ѝ���#Xs\PC3虼7=���r���;(�b8����9ϙ 䉣wэ��{U�M���K�P���=�M�9s׉@M�R�qR)f;Lj�j�'�M�7x�v%�*v�}���4��e��V#���O��^��A��	ו��p�P�]K\��R��W��
uC*�p��`E�AćoVyGW/ˮ*#Ҫ�(�v�*�O�S���}J�r�Va���������};�~5ʍ�Z^v[�k`�M��Z`"!|����9_?6)��DP�ntٞ��b��F�Ji��������8�qq)��#�I�ąq�*��-�-��K�y��ܬ���o�cl���E fh�B���cO�7���d�RL�ތ�6��'U��+���-'<W�Q���Z���`u[�|�w�t�Ʈ3'�k�l�[��L��1k�.]���/�G�}ls0�`�Ů���� ���?�7��ښ�1��O�W_�<N?��6 �	m�y�~��Pj�C���Չ���fKBZ�L�l��(#��
�PA�]�z�T�TGs�*nlkR��֮�X��e�/I�̜��|�:=�ߒk�5�|~4N'������k�u|�Uܹ�0l��[ۯ@2�^�L�n��Yc�:���ؖ����'[�v��~���S�i�)��Yy�j���"����y������C����/�B�D��v�k�⩝�G+�|�z~>�)h��~�^`��Yܫ���!�������^��4���或��08���ԑc��/�˘�ukm�j���S��1r����MygmM��\;�k��?i��>�^�v{)Ѣ`y���N͔�?V$�w��t��l������MO]�|u)e����V�����^c��U&w��q;ف�uiIvC���Oq���M���_��i<��{�9���)�����/k��?߻�HRRrg�/yzQ��t�U߃�z{�	�Ͼ��[��}�c@�0d������Eݏ-�X9��_�E�m<���z2�,X[Y��t�RK Vx2t7.9���y��\N�w'Ӱ.�j�>@�1�%�{t�q�a=o�V���;�]w��@WcL1c�qR�G�2ӃN��UE�ږ�����
IH�4f�$6K�v�������E��=�9�y���_�G�:Y�rbpO�u<�X:�>�[W����&� ���K�:ӂ��6e�}9��,[�����u��䧃����"�!ֵKOl.���l�D��}�I�T�O���2~����l�ڒ���P�#}�{�6$=�sPm�<��<}��q����5Kb�mwD�vM��[����%����?[�����7{�#mCS��;~�Zy`ıg���a؜po�*�/���]��%��7�7�����S}zQ�[�����1����fm��wa�� ����3���U]M��YQ���+mZ2K5^sw��-)��ְ�����S��G����e� ~UD��8����C��s����6����4�5��Z��G�Jt��d~�����y�̏�4h����CPS�&��j��ݍ=Nh�
{>w�݋u������Ǯ�a\::3���a�sd�"�d�*Ԁ��~��c��_����������
²����Z���~c��������ҁ�4��˴�}F�Z���KU;5[����5����%wdf�� Fot��{zD3��	��qx���J������*�M�����M�sh�����1r0��2ɻ��[��x�>���� /3 �k͛7a�`G�����6�@^L�)�ۡ.3�	tNkᯉ��H�A��0�-h:!_n�#��{��Y]�T���>�D�ɳ_�=&#�1Jʲ���^����gwO�� �'���׼���5��Į䢬��^9���`M�$���d�zpW����gűw�n��<I��l5}�s���O�:���������f^�j��z�r��<)Ҥ�l�!3����:��M<v�������3=�&U�j�!���\7�b�U8�����>ǘD}���1G/܈���Q�/��J8j��Hn��co�p6uwGn�@x�����d��J����M�°�޸ɚ���U~eI��*�'.y]��UԜ_�v���S��ߪ�����&^6��������؄�����Wbw����{���7���ձ��-L�r�v���n���?�6qu����~'��{�E���>���	5R�l<��)c����s	3@��շ�죇Zߵw����9�Ւ���CW���󅛗��B��L�"Q��9��Z�k���!�)�tJ�t���-�8��]�p���Z��&zS>➑�^��S���T���4��c�ŏ�a���f�9A��7-���K�e�~.�o(k��b=M�5�������/�6<�a�G��j��+�q��[_�5�,.�Y{bsf~����A����
f���ѭ�P�)������7���hu~�7�3c�n����s��I�6�NZ�2�^xгv��I�q{�����b��+�_px]����l�oS���*/j�i3��p�S��m�O	Y�~�I�XD߷����r��-l�+�b���,��g��1���Y3­���:�?>���t�����KC'OEgl�������$������n�S��6��+�v��E�W�4n�Q��Om�Eڍ�U���VE�kj����0i�͇��I����P�	;{;�y\P�(�ۑT(��c����MS�����W $uBPP�-�r���e��� �]:ć��~�~�]�4Wi��7���_�J�H�>����:5������?��آ}P�s���[_��s���ځg ��*�7'���C�'�>����=qΩ;s��+����3�Z�7�r��߭ĩ�ۗ�y���Sf���4�_q�B���9y�9J���k<gӤ#�{.NJO!w�o�~H�Wl��|A}��v�Y����g�*n4s(���L�˶s��xV�=y'��#�7�`sy�mJ��z݊h@9��v�5	9ő�_L�����ˋ�_H��Z���}R�1���lqi�h��a�!m]��j�ce��߸[��ـT_���v��{[-��F-y�O��[n�.^�>6'%@��W�g}��񋀱����=1��� Ӛ��R�V��uω{ݟ��*���V�m�GͶb�6�oX��.�r��ы��/?��w?���{;Z߃���z��W�#ߎ���}W���s�ܣ��Nw4�ѫ�^�1�_v��&���S�oB>�9S�c��k����*�X���Z~t�x+>����Q��7��T*5�����"�$u"1�u9���ƹ�pۢ�+RKj�P�a�-�뉻� ��.|�B������Х�ւwc������:��t�y|gu��`����i��c��Z�)O"���JY��I:(��|��H�����c~���Y��&�-���S1Ό>�CO5w��4��Q�h�͘��ރ�C��_���S8b��Uq���+�ʹ�O��a�3k��.���]`�+v�v��IN<�{��7Vi��ι^�Sg`ו�_��?;���n"�G{�vF�:��f����=�`����/=�U�lU����L�h�*k ~}>�L���7�u�Q�.�6�X��&�9�9P��t's�{�\PJ��[�|�=�\R��5�Ԣ��ƺ��+ϻ�VzjnZ|�o[��R-��'��/�ߔ_
XJ��|;�
Թ�T'c�W��nq���s����SQ0�zZ�ߋ���Pu�a_\����}�}֐/u!e��|�\�˕�n:/"�Uf��F=�!
��6�=���#�`�.���w	��_&��-y���&�5�ߗ�/'��5�����t�:�U�U�@5�5O[N :�*__*��^��A@dT�q�y�(�j��1o���M�j��ӎ�lڻ�;}��l�[if\^�)s��u{�a�=3�(ѓ����,�X[ЄUf�Fa��=� >{�".��K���-xr=�A����Fzƻ�即��f���=���x4�׫���ݧuo�ֆh:�l	��t�,����.�A��n܅�!Gg�'����(�prW%�Z�6��\��&TN��{��7����z�s�[}�Iz���f7ў�����^[�q�E�@|�I�٤]�nj��>�ч������Ќ�z�w~*�0���ȡߧzS>���S� �ʐG�ݛ?~������J����a��9
#DQ,��L\qg�q��gy���"���#.���Mlk�z<�y�����}��A�w�n�s4�۝����''.�����o>���p�k]T��뻓S��j�Cv}_�fe�5�A<���h�窋cΙX=3gG�}=��y�x��֫����??�C��������c!u�?�i�K�M�v�f|z��� ��dd2U�!���!��x���YO����~P��:���Z�����O��~�]-0��+ey���y��Io�Z������]���v���cm��o2Qڄ�����N���i5*��W]��8|z|l��->*��1|'chh>����徛2ރ��/?~��ĕ�n�����t��|�h�iq�L�q�inu���)�?tnN�
ϼ�{��������.��D�Fe7�,�r�B��++@f��������d\)-`ʸN\����A<�����������=�AW�nY~�W3�(��h��ŋ*^.���&��ߙ���Haɔb.�uB��d��k�_�eq|�,_��ˌ���9��7�k���T���j�@�1oh�V�7�jU��N/�U�k�Od�%̧S��a����8���F��b1?�sGK;�^�V���y��`t�L���^�/7Aw��
'�U�~i�6�F�M�Z|�)t�M��DZ�XF�t���&�b�xd��w���g��A�ߙ.;�f3`ٍMY��/��>�ܹ���\�Dj���\tTm��COD��}�*�N��:\�s���'>��MS��1Z�K�w��{�ˣ�j#�����~�q9t8�X�
�ӫ�����X��xmï
���N��^���խ�5h�{Ȥin�РS#��ի�hٖE)W�w6����i 0��o&b����$peLS��w39�Q���@�L����vL<|l����6��@1���w�r�a�vX �1���Aa���h�
� (�N�ۀ��,\���n���"�m ��A�Ap�G��\}+�]l�Z������bmk��`(ZY��YZ�YZ���0p\�pv�r��HN�L���n�Ll���Z�Z[��<�%����Y�+X$c*v��'�7�-�e|Q��_�3Y��n�5��r������y�!R�߳p�@��+�ɂ������ö�I�L�#S,��̿f�E��?s: ���?�	����݇]���=mP���&�`��@S�� ��0����y@���]g�\`�L$��D�?v�
!���>�l� ����;����q��] �.��l�,�m�@����?aD������+ƿ����X�[(���?�P�C�� &_��t��)������oӊ��`�_+u��,
����e�?f��fv�|���������˭�� .��/s��}�?n��F���8w����G����B&��� m�p"9�G��p
N�#�p�B�S1�r���B�N�nC�� ������71T���Ŀ/D8��;�YV8C�3�ȂcyDNE!xT4��A=p�P����"d���o@'����Gt�۸��P7'��F)(E(�f;+�~��E9#BٮNp���*	M���7����B%�����CQ�?"ñ$8�@Zg�-�3�/�(���iC�  `n_�)&*+,��Xfh����a�2Ct�ZK@P�ϴ0���U�(��-�$33[m�,����,ki�l�����%�����{t�qܰ�m��^(�T]�=(�U��?lt�+�����-!Nb�FT˷E�8�)#��Oh|�l���Ԫ��7��y�ؔ�e��ǳ�����ZA���'V{ܛ���Qq�NO��e<�n��EѢ�&���'�;�w#-�c�5OU:�}��ﮁF��-�o�pc�.�I�Z��b�]�����:r��K�����t�O��+s��]��Cn��* ���X�����,�?����wuX�L��V��	�ŝ�K����-��8$I�A���Ey/=�Ԭ&��ٻ�î�O�N����S��+�U開<�ύ	ӧ��Vc�����GQ����L�	U8=�hr({�	I���m�NN�OY0�����I���s�+$�#�X]/+A�RKQ�խH�u�V������������oP��iҖ�/=�A)"2Q�G�|�� 9)K��y�ܫ7Ȉw7BثC�߽�O��}<����6�s��}K�j�t_�
�sx�U\�䉢�oTBp������]T�A�MB���X��ݜ!e�)d
��k1D���A�y%] Q���>�Bf_�>#d2�J�p`"3i4]�r��kJ`E��dΏX�n��x�:�{��LL���"�G�k�Td�īw�Б�/P��ґB���t��?%
񾺀nd�I�b����ج �w�7��p��d��2%�0]��K\k_�I�
z��|{g�s��B@��	-/Gn�F�b���Wl`��P�R]m���@~�Rm��J:{|�������D�p�Z�5��s�]8����5 �CR�,�r+9�Z�J4��w��.K����/����4��<���U!�u*��բl	~/��t
�Ƨ}��^�o~�ɒLP�	!'2��!�\)p�l7M%�W6�u���-<e��/X�$�
9pIzp�~�����l�H09I
�5i�����&����6
ݸ��B����κD�3�X�ځ���\�*�	mV⑺�3A��m��k �u;�*N���󲿢���Y��,�'ԥlx=}�d�!��H�w��e{֔t'���Bρ
��[=0�^ �pw��i�
�����Oٴ� �v.J0�"8��ᭈ�Bɳ�͢Ȥ�e�y	�l1_�,�L�x�1��d,@p����u�
Vؔ�stj�;�l��h�cr6���&)�F�v��#bCo�"�)d�3-p���4Z�J�]h�\{V���Ƞ Jy������,��z�0<	b`���u#��6E�S�#>�'���ɲM&R��5|�2�~�Ԏ7�Ea�6����\P������U�d�0>�M�E�"hrB�i�P~�ɽ��Z��X^�Թ�8�,��J��R��j�}E�W�t2�8<mj��E�Ќ��<i*����dr���m�GfnoV��O|jυ������f�A��lr�W�Ϧ��3a�oT�f/��%��;������B�L$�V&Xk�GA�����ؤ�$�9�;À�����>-���~�{	��/�ɑqCC���R'�?*.:=��U�-̜'σ�8�y��SS[�U{mW�DtX%�Ka�%7�p���6ѓ�a�pQ������z�9�Izei�0���۸v�k�#u����3���H�3�l>+�e1�O5A���.oK,qewB�Xb*�����>@v&JQ�+mő��3cE�tt��<废���6���4�q-�QT;�jp��ߌ'�NQ�����=ɋ�w�|"��v��@�foٞ+xU~�qd����M;bS���Q;��qI���uԞ+d�T/�(�&ҹ�zٸYW�(y8u�7�2ƚe�3���G�Kj ��n�.M,���1�NS�
Zw��nq��P�ㅔ��,�Ւ��e�}�>pER8��O��UY��Az�ƹ�N	e|�J@���	�kP�'���%�/�Z9�KazoM+sʂ��p�҂��V��VK	0?hs�L�L;-p�/�;)��䰺���/D��bi�9�sV�#�mA��k|O��\/�u1���y�	W��5vO���u/D�µz~�o�����8����҈jz�V�$� �Hᨭ"D�"�5�@0/��+)[[�Q�(�[�������A�uw՜��:;�v����Z����4�0�Y	%�Ȫ��f�;Vwn��{��y"�fE[SU��F��pP� kO�g�g�+lSZ����;qɎ&R�CӠ�>�����H�n����f@1�����z���rU��6Q��It7����u�Y._����zb8�Lh~K;�Cw�TZZ$�3�q�g�<ZeӋ�<y:Y���/�����#�/d����V$��s�i�~�r��['vkq���`���!�V�R��ס1o��'����4uk<_�0����p�ۓ=�2/f3~��a���Z�=��׏�6�|x��SxD��-����t��q,v���*��J��Nq����:d)l�+�k�}�R=I:�� v��2`L[{��;����!��h��Y�PeX�0�b49�!���-҄<0V'
<�ꌶ�G"��+�e(H����\^�R�;�7 g�:ݺ<	�i�Vb�]|�O& ���Ro���F�i�j��PD�E>S�ɵ��P�1OHS�^�r�c�M8�|�g��W����X*����pl��Qd�eDH����H���|Pd����T�0�Fun����D�So[�c�i����r�ρ�YKB�����@�Ǉ���5�P@�	���|�h� >�V�d����ֻKw�-(^����M�MN�������D��S�Hv�j��E�W���>y������Z|ȋ8q�;R1��S��	�\_� �v�}�J�쇞���`m�S��:�O`Xl�H��'mi\�嘫6���"����ә�P�M$m����Y�B�wo.,�`C/8�\�,%Ɋ@I"��)�d�*�5Dq�@�~�����b��d�~2��QY�CxM��ǉrH��f�n(t��ܵz�b��/n���I 	~���H���?���c,�L��m ve?��HĻ�y�Q��,�A�vC�G����@c}]xHum �A�y�K L(%��zl�U�� O��F���kvڨ�|!_tT�}������d&���-(;�"�n��cSdDb�v��5��
�QeJH
9�������D����Ѥ	Ӭ�s9�`�^��Qx�
1𝈻�5j�e�[��S�H�����(﫬a6��LJ��ց�c�4ٙ?-�����������:��Ƙ�P��ƍ(�E�T�C[�p#=TK)E��ɺ'�,��Hl>;���*
YU�]�<p�F�L{�:����s��K�Q�����i���XU����d�U������g�D�u-ϟCZ�e��4�QGb���������gO1&9�Е@�8�<�u�g�8������;�'f��@PQ����e���q#�i�q�Q^k�V��
L�j�\	�	�}��HV�70���ن�H��C��љ�}~3^�ǁ��Ԉ���{:��T�L4�1@�����h[��(~fD�N����o����CX}o�y!�Q�H�!|M���������>���Mc�0�wh�\�1���r�+�t@.�u؅��� �E�R]������U<�T�c��i�n�
l�^��p�Kk1����'�o�;�m�e�qG$�횎% �E�,M�ORBj��R�i����v{�f�d{��T�$'�z��	���j8!'�A� �r�d�()X+Rc��?�mTr�ܱ�Dd 0K҆�(�?�69.֌͙kq�c��{���ͱ���Tv�s�bQ36>s�~�3����2l�6��8T�1Ճ��zO��5� �f�#�)c�چی��[U�å��	����		JL"2\�O�ު�`�ҍ�#y�xL٨2j`��J�y\@��F?m���\u>���]}9KQ��6�� �s�8�̝ʕw恂����n%�ב���퉥e�S�!�ʨ�-�N
[�)[�9&�c��4�6 �
Vmƅ=y �x��d�؏�"pۢ�:�9t��7��F������&,�Ԓ�v;��iy0�>�&Q�;~3'$���~>exc �g���d��o\�	)�덍-��O�}{���n`̝�-a�)^��u`�n5��sv\$�l�Yʉ��z�0	;�8��F>�8�ȱ�H_��s$u�u��� �ޱU�C}п���s��L�VuG;#c�@n�.&��mt��::U��U�E��>{ū54�B&l���iJ�iZ�Gw�Oo�\���HzaB��
�V��C7��V����e��)��zB�M��;��Z����'��s�N/�+N~�6�{B���L�Q����)�����N��CU���o$���_[md�pAe�G�\�X�Si9�"ŭh,���ι�d�n�<}z�$!�����:\nR�^�nan���8ڐ���Bdȱ���I�x�ɬ�!3>�z�:*�-��	P����L�nď��h}����H��D��ւ�(�K�U��cta�Az�Wy�^��f�ޛ��tňx��]��32������y���8u]?j�f ��9����٭�8�*��o�ݶm�dG�|T�F��	{T���Su%ˑ{���I�2��[(��.)���n�D`k�S|�!Q���O5��Lfbϕ`
���J���`�p08��7ea�,�~�8 ��>�߃�"
�" �2��Z��Hw%ר@��{�7V$9��Oe`��%��pf�-�\�yv�,�4�R(@t+��8P�Q�oH}r{�yS$TN� q�[L�I�|+})�,�D-,�
V�>}ÂL�C7S���aP���)5Jb �㻑���mAuQ�`}E[+T�y�s�w����;��X�j�-ܶs��J� O՞����iTxPO5�	�ӕGt�m���'�5�Y��d�$R!��o�okꋨvs�u[,i�x̌�J(d*�K�T{+?&�]涗�y��x;�)��X��gRY��׺���Q�߼�2><VH��mB?*���
���^��V��[Qcqu���#��s��O#EA�>Rդ4�j�l��O�̋^�y�S4j$�n:B!�$x�h����-������yK��,�}B�K��gv��e�/�Ѻ,(qY6# ﲤ�S8�mڿ_�@tJ��y��_t<��B�T�̋��@�pq�2����:� ��.��8B!�%.����^�:�4�>P���KG>E�	;
G���?�Po�Í���*�=���L�u�����+Q���Y����4³���e��v)[bnV���T�3ȴ�w���pO�疛-��HZ�S�5�\�_#�`r���@O���[_�3�8BV@)RRx4Xk$Ѕ�w'�0�纝i\�N֏
��/�X,����})�3m�.Io80�@)�1<���~�>��
S�G�5�w��?a����߿��j�uY�Q��T��B���<�
k��y��2+_Z`�@(��}����lث-������={̢?�y/����Ιw_�vp��p�c�S##�ݶ��/����T"�E�|a�zx1���ޓ�Yc�Y����Zۓ�?�~Y7}���zg���	�"�����v��It�w�~��|g����mJ�u�;��r1��]�3��p����d�z�j�<��J$��1��ֶ�Y���C��(���T�`����T���`-ZZnݳ(����	��C�7}�}�=κ(����-��+lu�f�����o#^?�j��|y��qtX|f�{4o��/,���} ��������@�A]W��OV��Ov7�:��#��o^|�R0��3����P����*���؝^�~6�kj}�?^�^���"�ić�D����Ϧe
���/ �z�F<C*�^h@@�I�d�B���хBz}8�N�O�Λ9��|[ֵ�Su�$���*M�$�ӻu� �$�s������T�%}N��V��\~�WV�^L��{5�w(���+�9�x/踍`�3�)��F���W�~JW.����%��׬6kĨ�_[f�Y`�� ��I��?N�T�/E���qjFBލ�õd��s�Dz*M�UQv�R�<��7��Qpt��������0H����s�s��k�*�AD�وE�������6�)�͏n��"�M����hzդ�`��@�(h��n���͑�_���+?N,�� <<����kl���:A�~��~-범��+p?�)��߲�rİwMe�2��^|Y�Qh���-ۏ�_)s��Z��������W�~���m��L�A���1W���G:�L���Y��3zM�>a�o�a�{5���ꍚŋ�������m_N�"yc��P��Wfsjӆ�0�0�:gu���3t/ҏ圈'�'z�����0FCo�=�G����?���T�S�u��ۿ���u�����{�����d�0�CmPo�F7)�*�QJ�~M��" y����z��S��.�p���߄���*������������7�pӯ/bI��F�b<ÑVE	 H�\5x�px�0�}3�c3�P{��#@U�\\U ���)A3�x�Y��H�P�95�˚(P{�$Gqt5 �H
������,�������do�${o<�9(��E�uY��H�!��Z�P<w��Q�0��'	�u���a�BKN��(�$�1B��@BpͱQ���%M���Hx7翕c)�����I�$�|H�fR�v���x����<�h�� �|UX4�� +���0$I�S�۾ya@P��$ꡕ�,A�]����5�[uH��ָ཮1c;.7/H��M2��
�q,�R�2$vZ�T]d�DD��:D 	WZi p)<  p4]u
���V5 �Hx��c<d��@����? ��� Sqs����� ���;]i�Խ����+x�x��+�/~�����dD�_h�8��+���Ѧ0/iO��`` ���_8���0Q��Ek�. ��;Qd!�����ía��eb -��glx���(�C�J�f��n��Wr��=��^ي�X�J��!���J�/3�.���x��UϹ?�xu�ya@0$�24OUܓ�⇚e��:���ၣJC5���[r	������в�}�<��0<\���G3]��"1�rQ���7�i����M�k^<�X�T�1��Њt�)�a<�swSo����Dp�{=�4���\3���6%8���jRK�G����IE�i��h1H�4�^;]'��45���e1@�TU� �8 Au�������ƾya@���$ CWܲb F�������r?�s�+�\������U�
�,�<X�|�#Sqڙ�8u�B+9�����t��G�ad&�\<h���WŕAT?��H���hF��Ga @�3���O�S#� 3ʯ�ԑ���� X��+*�\i�9o<C�ġ{A��h�@r$�VT)�F
)���Q��UJ4.\R�.���z7[ծ�A*`�?��.^d��I ��G|����<��0����W̰��n^�����Q<��Ŀ��O��#���������g��n�y�@ݘ��C`�\���W�H����!�ۡ�k�/����������#��K�C����ң�/�A�&��_BZ�ŮϽ���w��C��t�J]�0{�R���3��L>3���3��L>3yW����_��<n~�FΟ_v_�u��￡�Y����w�-�����qU~��﹑��W8��
�TP�i���|t��Z�H����p/�����/��_���*@��O�����cꎎ��>�l�A7�۷;%���ǟ_Nn=���e0���%_�����g�^�c�}����C]A
� `)��W$Ap8��$�ྖ���j8k��nT��ѯ;�"���QX�z8�y'�R��Gv@����ҵIU',�}�OR��)����-}�d8��C�%��u�k3�~�{�7�{���c̏=��䟥��^s����i�zT����.�����u	�$�c9�,?%�{�G2���}As_ƽ��Ɉ�q�/��z푄�/�5�C��׹�n�t�'�����о�(��F�׷'���~���ΰ)O���gӝ�����A���D�k
#AlBgU!���֑��)�v�_��VW�"�����4���w�L�>� �5Zh���EvBA�,pKh�����IS�&��dQ�u�;O=���n}���6D��v���aS��?�Du���,y�٭=����5[��V1C9�d�IZ|�v�|?��pT�P����kj�"mMP�*ZS0O�o	e�Ԧ���J®-�jiՅ*�����ԡPG�E�b��j�C��(���u�j	�����������ޔ�d3�g�I?�}qo��`(�N�������m3T��x��f԰�L�h����L�q�(��N���}o�wP�mF��+zWL4><�S�11�Rh`�LCޘ�~b���2�vFi��ڝ&�jj��gf+h��}P�q���#=L��z~����F��L��:a�d�)��d������U��:k�VYg~�!֛���)M4�o{�7oNc����-�)uI���y�4��監��fl�.RÑ�v��ޙ�vީȝ�\�g�H��������:׆G�3Z����ЙzbM%�N���NlIjɠ��׊Xk��a0_'�͙�j3X%�m��͆9�馶�MZ�$�Y"��^f4�6�r�PZ�,�'��/b��5�����!��͞S�N����<�Ms��>"D���n�-- 6����k=O�w�͏�?	#�Ix%��1��n��[�MsΤ�f$���N.YO�� ��t�9\��~'�~en�l�&f,�9	��^�+�YmM�J��K�~���*����a�wlݩyJ��a����w�k�֡��)�!�����m����<[��\+Ĳ.��9��E#���.���2�p�묡�ֺ�'������36�R�
�+�>s�gP]2��}b%�� mr��v���� ���n�T�����2��?i�&מ�37kq��q��h�r�A�
�*�iH,ƨ��L�ܫ���gl;t͎���Bۈ Ґ�2�m��lM����l������\��W8�V�=I�p}1�p{�05Z�'͈���|��Iig�)=��1k1[�a�����1~mZ# ��=*\�J�M�8 @�=w ��*�|w@�JG�b�o=�J��p�d�X#�$p�u�b�u^Ѭ��o�k��E���oj+��3�M�6�Ƚ���{�1��M#���Ѡ��Z�p�:	�M�ް�hv�E\#a�Vh��q1e��Ƒ5
��ӈGٲ�������5�z�N�(�ǵ����I�TC1's��S�aE����\�Q����(T���nm�������찓�!o���1Ӡ���~v>F71<Sj�S�5��!�@��� �jĔV�6�qLz�x�G%�P#G�i�Ӗ�q�V���^"����C�@��υ6m�V���wm����T��|,
"j���b6q�邭���g�l�Ԏ�^Ϸ=���eq&����i�H�36�v�[�qEm
z���#�'v�rؕ�H9��8Ms=D���;P���x�v�;o.�N�=[6gt���r��L�Tu�q>�C�D���"m�� ���N�t㒾C��Y`/��YI[�Z:j�%Z%��f�4��� �;��T�A*vn]Y������3�\�kTX�H�Cb��� ��dȬl�ZbkCutF ��k�]�'k]���ͦ��IA`V�4)�w�w)�%��4�L�ok�,�R�G-M,;sz;-��(v�d�X�{��4GYźgȚC���t���^:�l�̭��i)t�㍭�$9
��C?�`�hh��J�XS�[��9]�#�m��JhX[�Mύ2��#��8�ѦYg.�K~r��)�ӧ974�A��G-WZ��ZS@v��,w{A�L�m?O��Hue؊��-i��������u/��#��Dl?x��j�h'کuO �[�4���I sP�����w����lL�[�V7ƥ�l�>�g\{8�B���TM%�ֵ�}����I��y��N���zݍU�M�U�DB=���&�b�i�g�4�)a�����=#�hDB�m��7����u�����p;By���n_6|��Izo��؈���������h��/gP	��N�`�L�c�=	�Y%n���V]��*QpAH*2$Hj� M��$5Qd����7PN�
�Կ��n��Y�M>�kDy����@�}�9���Be�yg�Żv  �ZI���z=@�9!�u1�D�HBw�����_+�o쀹
��Ƈ1~X ޫ�;��rSz����|�M�`Q������(�N�BOK����]��a�W�˓�����	��jQ�H�ɨ�a���DB�f1{�,~�?:w󭝼:>����w:�于�ծg�88 �V����?����>��rv<l���uBT.���-p�wY=�	Mo�#r�����Nd����"bW�;���w5��(���l����V������)�����#y�n0{�*�0cZ�j;'/-y����)������R~ėl�O�p4�)�ӆ�4.$��8'���u�u-`"M�^ؗ����S���s�=��I��&�C�kՑ�@~�H��|O،4L��~By�bW�YN�=^�+3�C�#"�Ƽ~���Yo�q��wx2�Y�AW����F�b��>ė0��g�8� �O)�����f�y��oSڽX¶�:?�(�+�:�5aϛ(�g	�O�
R�m�+$��$Iйs���|JdcV����V������	T�9�.����P@�)��_C�'����q���9a^΢O+̜35���?��!	�Oͨ�_mu|�#sϐ)t��A�a�d���<}��BI�a��m��K�Z�䗾tw����p�4��	��j�ۘ�q��qN�]w��d0|.�u)�q�TR�m�VF{4�x��09ea4���@����5�NC�^M_�E3���+g)o���X��|�Zrb�~�8�~�s��T/��#�����L�p,u�`����P�OG�g��C����!$�㓕+Q�����S�)onAK���㖆7���zi`�$���{��m��GC�Q9�3��Ni��d��]���T8�7.���%t�>{�rq�����!��5Җ�?#���<�
����6�Ͽl�s�C�8h���QSW>��3Y�e`h��%\#:�7�^��˗�N�<O�C��_�	�?�p/�1��D=��s_�`m���t��Y=n>�<�<O ��Q5�#FH(A�_�Sc�n�6޽/�t�DD���ɶ��x��l:%�K#e�(0e�uu?�E���> %��)�\XQ��v^39��(���Q4��Z痗��Vfu�&�>l���U�Yw=d���h����$�)O�<{ܯ�l#�қ�H�^�;\x�h'մ����R�q�6�~�7�@I�R�K�)�6OS��.A��_@CM��6u/�u�-�?\ƺ��`�Y���Hn��U�B|� 7�ph忟�Tnxt���6����x�^ �CK�]ɒ�Hr��2�#m�}����$@� ��"@�ľ� ��]t�i���H��P0�Ykf-�nu�H�f�$�၈��y���a/A���Ɂ�c �ق�0<������B�@��[�:��|&�Ѷ�1�I�|EF&��9���f�(_��Ợ��_�P �>@F����sU��Rt�c!��r�#q���Sw]f�	��򓦠dG,�݀y5v�v�\̽t�Q���Qg��!����*�A$��(�W�Մ6]M�D߮�>��#CL��nS������ێ0*A ��C<�ry��V�֘A������"kO@��:ɮ�T��"� �v4�|���+1.�i�|~T�s�2K�_�z�R=��G��$�����тܢQ��'�좎[U�� �V#^38��dX_�WI��D9\����Ȫ���6{NaV9ۅL<Wc�����p�do��#pVZѓ
�1^Y��ZW�����O���^�xwQ4�Z�+5H���l�Z-����3�]F�3n��v��=,U��yd��̵$��'��(ahÜX����Ђ~ࣇ,Ef#VC����氉��bh�8b��J<�$t�})���|p�V�)�
�j��hB����CeTW[��b�PDR�j���8���Nד`O{���v�DK �2T.��1�HME��e�\��X�< ��q�� @��>�R�%
{'�k�x�C�����I;T!�2,�0tX+��t�ԚZH>[��|�m�"����ȅ�-���$0���IR_��ԉf�����:� �0z������Vv'�i�A��5\wO*��d�,s��Qw^E3_�^U���`𓖈4M�5�� eBQ�Velh����CT�ઇ8�N�=��CT��S	؄	�=p���gX�E	5�aP־ݴs%Q�Z� ʰ��Q��$�x+�����^�R����^�U����&Y�Q�z�ꊕ\%p=G26n�!��u��Ӹ�G@�z��u������I������A/�����u���E8X|/`|dQ�~�x��F=�`�lt)BXK���GI8`�-�D|S����D�`r��7�2:��n��U�菆����p�*��ݶv��^ʜ�c���ӽ��3Y�-c�#D�2��,�BW�.���dXi�{�%ZI�r�;�nUK߯���B����=���ILi���.��`��ËF�t��C.��m����g�(W��#6B$�^���ř��ō ��ø> v&�X�=_�Y�d�vێ`)I�����7�v��#�\�]g��̄�>�nw���K"R��Ʋbt0 ~�Y��s�+:�s��$�^\�+�ų=��*�-@�{ �~ǰ�yW��M:+̖)��ŚMu���������,2b���1(z[��aj�d\]�������g��XDN��:��^�c��j�_.W2�&ԧ���K�A%{�[)�#�a}Q��f�a�	���kS�����E�UY��yG����&P�}���w�'�B�τ��';5=\�
�d���ٵ��!38����i~1A���N�ti��\V�t9����<�w�[kR�,�o��P���s9@�|+�uvJ$=u��`Ռ�3��9G�vs�$o�W�f�.Ǎ��k*�h(b�Ս���J���.�'��.QVn�4]�i�.��0i3�!S,�b,W����@�8�bҦ]u^&�Nb&ˠ糁+̲x�`�cZ�.���.@|��ˆ�Pa�Z��q�̺��8��`������vL����e�� T�4�[�<���Vm��dĄmJ�b�lAȎdr:�p�21�'�#͆M �8l,O��r�-�"��
qE¦d,�J���F�VC�ƫ����aB�Q5FR	}&g�ڻ��l���$7P��S��n���>h��>�
����V�_�ḛH.��d1n�M�V�~��[;�K�M�l��R7�:Ԓ� �h~�^o5����G[�ZW��r��^��eKE�T����)c��z����Α�*:�B�����3�K ݛ���U]!.qC���u�ٯ�qgI�urW����Eۋ�bg^ņ�Qg�`�9xx� U��L�=?䱺��Zh�o,�1���:���9�u�ԱU��NR�2;|0�}
0�v����E��M�KD2��Y�!�NtB���!�<|�Ǟ��Yj�E�o���EMW�vKwR\t?�����{�J|=rKgRJ�U�;8����ō������N�I����XǄ����u�ل?e\3˥��V�!ﱰ,(:��X��T�r��,�IR[1�@������'-SO(��o���a��_yg���'u)���Q���t�zx������,!������үn�A�ٽ��K�����Qd�괽\��%�NZ�3�TºFO�B�pe��Q�a[��V,`��q�s�T~1�O��<i�%�{��/�I�"���'KM���&Z�\�]l�Ę�,B�R�%Z;�)�2�mNY�p�4�fl�^'S՚6��n���N"YhT�2"[��0��Z����JWs�V�?���!��5�YU�d��)��s4GD3j�ĩ��+��aͲ����>�<��������$yM;B�E�]�l��ᰙȭDDt���P�I�j��]9l����Y}�i�� �g�3K�vG{�w��E�M*�6����`~��������3uЪ�:��A{d�����r ��3���Վ:P!�4u>če��&�F^��`H�{C������P����=��ȼG�_zQ�9yd�G��u{�nV
J����m	��í^��mz���bfE&X�S�lZW�
s����L�䡡��� R4������0+�;JK`�C�I��}^Ƙt�=I����i.�����J��唣,{1]�iwA���c��s ��ˌ���FB��>́R0�:ꃃX�7����qo��i�����4���ۙ@�8)`I�� ,/���a�i�V�鳦/q>~wKP{�|��4}�sQG�(wS�=Y��,0�	Ks<� ��,�(C�$����_h���}<��O���YCa!*Ƴ�l˱��~:9�㦟���S��l_�xo5mQ_^�{�]����%���?*�_�}P��B]�!��͂6����&�/�-�i������Ic��)r�}~��ی�o2���c�w*�'M_�>�S&"�g��-��ő�L��^g�a{v뀽�x�ZJ�K����On~�s����+�XH�_?��ϯ������l�T?_}'�E_��6w;�W���QS����B����Gٷ`=@�x���(�߄��_ɶ�Z�����6��*����|;��y{�_������N�����K/vy�>,s�4τ��^x���~aH�۽�yG�t�sʅ�Qyi��nހ��yݴ	޵~��K�6����5l��^����s6�%~)��+�	��m��T	�>h�y���Gw��Xt�(��������c]�.������o�|�}�A>l�����SK0�7ܷ`����$��|�u&@��o���YJ>���1Gi0κ�Ϗ?SU����o�Gs�L�{{ӏ����(�.?�ž=���5�v�]����_��_��0�SJ��M�on�-#����MR�_����w���)F���IP��4�<dJM���0yzyͦ���xy�wit�����������	�.8v�[�e[���M$���%�۴O���0^�����g�z�g��n��I�}���Ϳ&��X,�t�EɾB�x��e8^�_�P���ءy�.r�u�|�]ھ����S	��D_��(����^����6��x��<��*������_����DU׉)��}g	8��2$�+�T0�"}�,0�!q ?�9�~�?Q�ujJ!4|�ap$<�����G2S%�w%��SpjJb(A�����k���X
��{ϝ&�)�(B�-���>��>`(��\�����!�aG��0L�w��LQ�D�Q`@b�N����)NP��E~����"����La��;���$��,���1�����B���gr����;����@N)��&pt��(F�C�疝�Gy��1eP
#�j�@�����q�H�B��AQ��;��4b ��)x˧��7�*UQ/*UJ��/�Uq�H���B�����ٚKX�{��﫟p;�Up@'��(;���'�Ah" ���4o���rܾڎ��I����"IP���@x���$��UI	7�L
�H��A��u����ɠ��"ԋI���D`�J!Pψ�ݎ���Y��T���漏�Ң����uU�˟5��F"��B|/�a���h�CqY�;��zV/D����i9Dah������8���:je>�1�ċaމ��f5ݮ����(�̵��#�a�7��:˿��Z>�d�}���ɔS���rZ���b#�tY��\;KTt ����<��7���/m��K�!0)�!x��Y�f�9�.Z{e1X�i��nZI#"�5��Gx���hϮM��	����*��@u_�ժ��qQ�h�@�A'���{�.�.R9� y��P���}mv^�^�#��e��1��!{��0>5��V���%� ��xh<�{9��匾f_8i����{;�4=�9��|j�T<T&ą�29��8�L0�����j��C")�}�֪0'���{�CF�{��U-D��B��h��qdtJ��p,�X�MSW�͈��e#+��1bb��U�`R97�P�n���b6e
m�̐�"Rp��U)i_}[Mf� �%h������@!����cA�i_|�&*Q�|kL�6R�Cˀ�c3 �v\5�sd��_w�g��hm��</�b�p�R|��TQ��P|ŧ@�vrю`���>=��-}�H�ա�LX \���?��!�uV{H S�����W&��Vx})c��٭�����|���;���OO|�{�E�"e��HYD�"�y���t �CK��u\To�>
ۍ݁��N�Nw�0�ݣ����b*��X���b�� �v��;�������������|�Ŭ�����Xk}�����/5�'*�k@�3DeVF�y�bc���~;�v���e��ШPȟQQ@�� O@��Qx�" ��g����6� �!p��� ��z����>��L�Ch�o�[�l�کW7��&O������Tz�ж:�'��a��6����-	���:ϥ���gd�q]F<��+�;]φ8�=�%Y=�u���M�դS��N?�$۾[|��l����ySª��Y�hې!�%�q�x�5uϴ�{�	��J���P��0!"z�natUM�׸��s�.8�����ô�)GNܻ8�
A�{������7��vpb�MSN8����/�B��a�}��t	J�m����=a��߷��_�1sπ�����֒�_�����?g�}[�������^�>>��$�=��k��-z�y�����'��4��_DLP'�̺���˃6����z���:~��K�@;��~8���}�bC�ӊ=�*ۆ<t��I������1ލ����|nh��=��-��� -CU�Ļ���g�v�i��S���G���c�f��1��qC�h��s�8��@펐 �s��[�X�w6������?�\��-�s�O)�DC��^S����ȿ��ſ���e^@EUvx���PL��u�x�?I̢�����[����A�S�ϫ�T�āB���"�p`�w��{����(�_;��CP;�@)(�����i�m��y!�l O�U^��?��*�S�w(0W��ҁ�\˟n��:����bb�5�3�6�,��� �aS䕙"Ӫ����o�v��{"�o��r4;��/���u����1�k-�~��ɟO�9P�!���}y%�r�o����HGzb�o�Z�x��}�o��4�>���-���[[~�Ȩ[&������t�1v������s�㿊jdm�*�>����}��Y����_?-�8��gۗ6�o���nIn��H�u���E����؇n��~x�:�W}h����k���+4�#p|������觸��_�?�����q�������t�����e�M=
?��xJ���ݶ漚OZ�#��M��NM��=�-�(��y���pk�L�Ş��y4f���~�9�ϟ.R�b�5�h��O���"�hr��۲w�m��3�ض>�m̇ܘ�[y}hyc��P��qO<�?���m?�������AA]��S�-H��}M؜�u3�r]�O���U�_0�>����'$�d�O;t୛nx��O��Y�vc�v���N���ɘ�e�&1kY˜�a�t�߱��t�s�p1�$?O�8�A���U��}�pA���Rt;:zs�����S1��������#W����Zb�${������>�w�=���C%��c\-�z�����E��<9�S�y�L��)E((����J��6����E�6�r��w�{ͺ=Ȱ��V�n-��V�*����ՖTW�6�R�T�J��4P��I����yE7�\5`���ﯼ����[ԯ�y7ծ^Y���E	���ޝ	V9�rVX��Q���q�ӵϥA(	A�q�1��[�*+1}����i�W����Z>>�����}�ƹ�}A��o�.���l�I_z����������T�%~�t�uR��CC��g���Q4����|��b�B���5�#��r�o���q�?"^É_��mAD	rF	�v��]���:sXf�����N��]���e"z�����{#����uU��r�MI�"�۴�T���=�D~�y�f��7����6�y=td��ea�����8o�*�����krSߘ`�ٛO/�r�~�^]m0f�Y�׻��b�6�e{�6��JD�r�'��޹ӭ�������v��o��Q�4�,!|S�fm:�[v�O�:���A`y��j��r�L�Ո�/�&q�9v_�qb��̔�?���յ5��%�{X�cg(�Hk���q�[��o[D����? 4�h �'Ԟ>�j����@�Y�/������`��6j�2EL����VrL��h�����T->�9ܮ��ux�iH�ñ{�.Q��d����$6�"%4	~�s��1��;�\���E�ط��"�2���=��es/�L7��J]v�'����+p\���z���U�<i}����S���K:ݨ%>N7}�|��sѶ�o7~b5��z���x���m�0t���Zp���h=wd�����ɨڍ�+�va\��sx{5���N���o���<K �@MK�K����5� l��3k��-���QU������w���Z�3{_�f\,wR�eX[�^_c%$˓.xM��/c���4gף	�;k_~�EF�o��t��]?f`��'��vG��Q�M�wK�ꟼq�f��f�u*h�V��	�ѳ���d�d��I�����-Ƨ��^�����j�z�`q^�G�#���[��t���J��ǟ��$m����b[ճ���6��\����꠲�]��j<A�'��y��߭����T�rJ���:�e֤���k�4.���g����s�_e��D�B���`4=�ɑY
e���d��^Et��K|O^v:��p�ǆk��G6w�wⷴ1S4��U�;~�����+T�0��dՎ�/>����;2)��es�ڑ�m�d���I��U�}���3�-�N��q�xS��S�MA�*��	"����ݠ=����d��W��H>w�,�z(z]`�nt�q6��0~z�U�����C�w�}�׽7i��|M���o�?��f�"���»-��&~,,���P�Y{�΢��~�;���^)/yG.*�;���RA9��U�g}�FTǠ�6��X��m胻uY��NW�G',�r~N����6^zN�����<xm�絑#��s�^�s�<�JT�e�!w^��ހ#�O�/��\�Z����{�{��Q���<`X�zڞ/n�f�̪�nc����tyf��>Ƌ�=4�a�;���kz,�:��j��Snv���௯(Jꍈ��y�(m�Ŷ�ϧ�0++E]�+];~,/{>fAj�E={-?S��+�~�f��C�{l`��W<��3s�,�Lm��&ݤi =SV`G.�ĥ��]����lB?lȥ�/"�/s2���T"��U
���H�ǽ�����.YG��yN�<�Z�����ߍ/�j�B�Jx<�-&��e��h�=r�d"�MѺ�aۓ��&���aZ��K�7���3f`&��(>aҘ��I��\�s=�X�u\��u2-�W�f�u��==}󸔡����d�Q�����
LH�->0�9�Ã���7�Sʭb����+>=,�5g���.�o�}�� ~g.}���J�����ۙN�����������gɡ�A7����
�م��3�����C۶���K��NbT�I7�����F�VVȪ��.��>x�"g�$4�P�-r�=`�������rT�؏K���A�Z��G'=�F�g*��hz�;l-a��Ү��=�}G��q�ݳ���x׍	�����⾑;�{��	-��,�X��n���^q?
���|�NZ6�1��#�X;���̹����o�8�l`�#C���a�?�� ��^�tb��S��M �ZxWh/k���/�+�}�6<�唺=����=d���oJz?�}����f�Ac_��o�r�%��ca��{�-�_���h�t�ɕG��/m���S:*4�s
�z�s�8��S'���Ϭ�	[p1(�'ׁ�\\ۋ���%���F�$�QG.��M�fX7h�L���Mط�;��Ӟ���n۽l�w��I�o��6�|\>��[���(U�v�kHfɓ)�EDM���Z��������딒�O/2e�
�a��SۗN�ߛ�d�Ҭ̛[�	�q����ZK���O��$���}���(��nje"�s�����k���˜�1CH�;�ރ>}����
�<�ȭ�|:�he��v�����`�L���hX����z�^b(m�?�_��������K� �w�􊶍k.>���ng�3Jo�}t�9�j��΃���x'O��F�H�/�ws�܉Mz)S~���D��'&��n+��7�lMn�p����|i��&?�.�؃}a�K� jKj�ak����k�o��nJ���;��}��t\�ݕ<z���ބ) �`��[�ujs�>��~�����Y����h�Ҡ/߃��e�C�ؗ\��^y�(>+u���InиX���!3b��6,��IM;�2���g¶��uY���V��.�7-f�Ӽ�>X�����3프��mz���9�z��i.���.ڟ0�K4o�8�O��wt�_��~�K�>�k؅�o�Y�E�����"�{g�'ƞ[�	)f��>������c���6'hJ/M��y���~r����N��-�@�|�7�}+�]9[�ר>��.�'�+ؑβ�Ǯ����ZT<�Xꑣ�v,�:+���"߷�����mx���r�&��կVr�]�W
���ӕ����;äjVQ��v�=r���;��vl^�����q���u�Ƹ^|۟:�NqE�"�S�x��6hW��c\co��ym�Z�I��iD���Ĝ����ͼ����}1�祷-���5��ؕˏ��-��i��D[��gjbS����4�k� 
�y}�ԙ�'[%�׳�3���_<ܿ��M�#a�M�ƈ;h��C��
��A�.{������.A��yA�H�sv��@K]S\̻��]#]��/&�K�����]�[����� ï$V�A�����U�h�L�_�{���=�{ᷖ��o�-HМ�i+y�~��+OD�s�-l����mt���?6�n�7��یS��}�GM�����c��ļokO�8�z=0&4��=a���f���9P��++{�b���}#�=(Z����hƕ��y�^�B�M۵�llT�o{s9ߺbמ�9w|�Q��E��[^�G_蒴�x�o����r�J��IV��7�?$���⽣h�6Ƕ?w��%g�D6f��ss���݆TL��ht�<4�׋/C���^�8gYy�ԝ7F��k���^�(��f��z/���.���?�	�,��[����	����s���O���N��=��,m��V䱇)B����J��W�0b6?�9qՠ�ui6ZkO�Z����OZl��(�7����;��j?|r�u�$bgJƷ�;wk���+#��G�:w�ҷ�Pɠ�����O�oW.�S�5�>	��P�c0�����Ҏ�21zj�s���?�>�b]N���*ָ�Jp]���U-~�LX&�!��|vL� �w�͸7�� qZXF��z��	��_�K��5aZ�/ī�1���pv�;?t]˽bD�1ُ��
|U��j����C;�?xp�bY��x���+6:�K#�v*���1�L	뗯^3=QX����w����6{��g���*���Boʼ�ƞ�~�~��
�yiD�C����]�9�ɜ�}��3=�i�0t�ZD��c˿�w!��`����j�@�1b�{e����Zql9p�~>�3�R�yW�Z}2y��O9��f6�d����Lg�m𡣫�����9���o�,R0;����P�Ê����E���.��ڽ]�-�~_�������z����KxH�X�%T�<�8�]?\���!��p=�;54�"���;���S�6c����<�t�m�a3�U_{M�t��8rб���7�:�e�n	7mr�,���C���Ǟ���r{�7���C^2��X�N���x��P����}O��MG�E����9|�t]bi8�`�y[`Ϋ1K���2��0����U�Y��3!��=sjǙ�ߵ����i�y��16��\���rb���Ե��/L�X�^���B���=�Ӆ�EG��o�-�q{�7�Ȯ����Q+�/T�ߴ�����h��k�C��˃*|���qa���nصt��jY����%���R���hU�l0�B����A�t�<x)�R7��L����ܽ��� 7r��[oM���T�#o�U4{��c�����spį�c"����Ƕ�����s���r}���w�w����2m�Z8� �p�7���ɳ���,/#����io�����e���*h,�Z[�<h�a���R4��Q>eG��9�vF�?u{32�x�k����4	%]\�Ol^Kk�3t�DLv��~��gR���IB�3�ކ��-	k��~���C�Ö�!���t8���1���e�3���C��+$to�<��Yp�����ۆ>���,|e�v��$3����?;ݥ(>j�w=iVY/-��8�6Go&��#1��=Ь==��F|~�+��=s��x`-��'m:�������� ��'֏)N_���2d������w춢�vU�}��&nd�����L�wr����6?��2���8R�T��vx8�i��nr�v沋�����ݴ��ۆ1��[��ލ۔S܎������_�[�IV�����uV�S��e6��Q�/�8�6��V�8��IFԕM1A�~��W�s*�)��J�f�����e�t�U��-;G]Qn{�c@���	;�_�!�N��V3N9	������C���ˎ,�{�/���,��T�U��ƌ=��p��J�Q׮�Y�>�l�
,���:i�-��p�=^��k~,�31j���sv-�t{�-�C懩e�&�vv&�ӎ��̞U[�<y���Y���t}N�����J��<��+[#ߙbﬁ���_��L~]�~���o? ��~m=T��}�b��J`/@k�|b�{���2ﯡ�Gu7X��U_�^���іҽk�_!��w�w;�BJg��w=����.��J�z_�<��y ��K���k�̥֒�Ϥ�1tK�<qOx������{~j�4CncӴ������$��_�G�\�(Z��}����(yУ�tPzn���Q����ei%��\��W�����\�ԅ�j�m��򏡋[^nu&��ׁ_�Y�Q�6��)����s�l���T�<TW窯�?���[?���-�ȩ!��kVu��m�ކ�N6J�<;�iBh���Z����������(���A�&�tݥ�U���ի������V����5$nؤ=�}��n�����L�_�Q;w�ް�����¨��e�ǳ���%_b�O�\�A��^wpReU��U�2����.5�nѓ�����nM�8yڊ�y���Έ!]G�6��q��{m�����"�����k��V���_68k���>�9���a�TL��)�{'��/;�{���g�[^nH{<>k���e�ԧk���A�2���Hޱ�H��������{��w���b{�m�r��R�n:�f��}i����So����۸�)��i[��\������|� ���oeͭ�7�V�"��GEߔ�4��ۡM����&�m����{	$Ҡ<��y�V�?%�cfw�`�7�Cy��7`Ӛ�BFÔk+J���=՝Wlx2t���U�[�d�n_�ܸ�y�./���$�{��1���dY�C��k�F1�Tl�� r�>�6�꭮�
���������^|T~��b�S��K�U/=w�s�����Ԍ����,3÷��񡫕<�y��En�'��Q��g�[�W<,���[)���1�bg����]&"�u+�,��cv��1�Β�}m�F(~+�G+�ʌ7�o
_��aIz���/�fY�C�"#�������ְa���
䆞oY����٥�����Mf�g-{$�.�n=�m�q�는ލI�IK����DՑ(|/��-q�*g��s����I�kmf��=!���2�|ԐO�-���F�e��p#�?�+ȑ����~��G��?����|<j`��_�f2�ա9��gwGJ#���\2R��oa[C��3�����b�N;�w�\Ex�#�7#l�5~�Ȥ;������BY���d���E،̤��?C^v?R�,<x���֗��B��.���`:[7�B�]�-ݑ��+>a���M��M�m���\	{v����%���o����������l�듇̃$��ܻ,��`7�bX�|�hrФ#�>�MM����z��~5���N��=�׬��[�̄�8��{�6��KfN}��tu n�4�����{��K�r@\o���=v|�nGk�3�͐}���d����ҽ���G����:��G���yS41-u�r������ګ{�a�85���h��}:����_=��)�_4������'�|�(sf��{��:�}Y�7l�g^���O]]�uZ����ؐ�h[��O{���2[�\�l�=���g5�n��s�3�|Iy5���h�g�������G���tU�>�x�$�-$xQ=�oO�~=����G��J�fX@���8�<z��'_T���"��%훸ԴR��F�u_��&y�U~�"����֙&��՞��_(]�T�'ŷ˲Ǝt�Y��X{�I%lK��>jM���~�S�}э�7�XF#�TS<�{��}Bs?}XҾ��λ�q7"d?v9G�Ls|�Sݫ��m2�ZP��cTY�#��F|��Я��GhVd���E96_�ž�|%��'���l�v-D�z���x������OF�8 ~�_��p�o��o[�Y�s�4:�f�J˳���.)��t�e]�O���ISk�90�c�TTp��#���R�z�ִ<�y>n��z��֒��u߀��{�[��ύ��G�]A��ƦUM�K��_�
�x�{�P��\"���|9��S�~�[��ܼ�w	.cl��U/�|���|_t��]��Q�9�WO?�����[z��`�Յ���ؠzN��9�3oɏ}N���|ц�ٽn"�Ʀ�� ?KI�\t��s�1��v�zr�>"�ғa���#C/{)��-�1q� n��Hݝ!���*��Pf�G<|n⪄��5�x�j,������tl-?�ۆ�W�ߞ�s��*௢/+��Fi�H9*Έ��Uب�+X��;��cp�H���a�_w�Nѩ��X����B����ϺO+4��ənI(g�@��@��X~}%j*wjY�8�Stص�G�'�q/�v��s�Έ�z�Y�ץ������.�}�Q���k�����ӤS��RsZ2޾��~�)����ߏ���Z��}��U;�a�{AɝS�=�gFP-���sRnV��yۿ�GuIW��ǋ�e��������\I�4=��r:�yT��� s��Щ�Tܔ5��Իf�"�n<�:&�-���U�̮��ȩ�K�^����d�β�Q�����]��-�]ݽ�oKP��wH�O[�I[���ٵ����&ч�.��Y�~�Q��7'�3c1�z��ah(=n���3������a"�����#�N�#�$Y�dN�s�w�՜�������>h������V�N&=-�,�k�TS}���|�)�Eґ3/?F��[>�v�5��lXr���k~٤<��ݚH���ݔ��=g0��uw�tgI�'ȟ����)'�b}l����GiO�*�z'�	6���O��av$��ݎ�]��G�=��)�A[jf����(����ʮ>��#.�2���U�^�Ӷ��G��$�я�+ח-�ڹ�l9�-ݓ�j<;7c�}h4�rM��./�ݟ��h]c_��!O
��W�+�#�mw��~/+�}�zzF{���QU�C7�Z��|�boq�1���gr��P�m�W���0������Ä�1�K��Zd��.��������ȯ�\��|e�04:tbދ��s�bn���u��ڰs%�M����ӃyhՉ5m�ff֙��JX��h�ۉ�� K�v��/6=�{�7�k�����/{×#�%7���:3��+�¼��>�&X�߳�@���`��M[�|^���)�gu���/ڣ����(�uD�8��ăj��7'��y�Xݚ3��X�(kTׯ���b~O9����IJGUs�?������hԆ��yA��qA�G�|�(���Pl��[a��7��ߵ�����o�?/^r3}��3�d������r Q����wەʪ��K��Z�q�|���Q�G��z5���8R������od6J
���r� ��Hs���l�-1s�]ߜ�H~g��:�K�����صܳS '��V�8m���uİ��-k��.��niZ���e�����`Ŝ�����ۗ��x�\�ʄ��k���'�~9rLE�f��#��0g���}?�l����v2�v�S��QU 6'�ę���Ȗ}��/O5�w�<��g�b1����9�v�c?B�ފ锶���^7g9#9�?��`<��'���y��@�1�y������NAC��:i�����+�D���1�P>���Q}��*��}�ا��Nͽ��h�������ڴm�Ⱊ������5�S�F.[�\����q�ſ����x��O�Sx����Ls����M��%ov=�u6��6���F�sj\w܃��\�����8����]���]~dzȂ��f���TvTF�r��>k�"�+��L�u>�V�k��u!=��,YBCI��FN���2�ͭ����Ǳ�-���J��HBo�y#���Ps���O�Q��#��H��R���`�t&�Q��gLnd�E���Qllڦ���u�0��t�ƁU7�J��7���E����-*{X ���p�e��1�G�.�E3��~gz.���)�X�0c{�:��0�����Ʒi�{J��4��z�`�h�P[���1֥�^焑��GC�/���땂�WS�X�K_Dt��^��_E��o�>ꤹ�~��S�)���Y^���'�~m��������������HY��g�M���4�n'��5,�@���qoi\�[sn<ۗwm'����"$g�9\tg��W��7 Z}��߂��}����6l�'��(���ּ��?�d�Q/^��$�xF�q�ɬi,=-?�H�a/��^T�\|����CL�M;�Q{g֌ޣ�3E�kQ�Gp�nN����?�V֍��oo����4Ԅ��P�����_�^���=h3�V1P�̙p,���q0o��߮s���yqN2j��V�C�'g�ۚbELfL�����ܥkS7I�������s��ӫ��e��.(3������hp��[����tG�[KQK�� VY���Py�i{��I���ھ���U�=vt�Π֝��W�z*?'pc�\�ڸ5d����=6��*�,���F`v6,��e�;C>w���\���܏o�2�[7�ڕ���ْQvtz�^/��6�C�ŉ�xU���֒�k��p�o[@e��خ�đ��x!/��_�5��JVy��{_��ͷK��N�pm�pw�f��9��.]8�j�oK%���Jq����]�jf5����eQ媢	��zEe��ݯV�7��b�����6@RRn��N��=Xvn��<`Fծ��8��sx�����]XF�_�Y���/��(���P��R˾�7_mo�/�7�؛v�L�nxQ�mە(���'oR��q���=�:-��h�.,ir��qٜl��!����^��V3�ki��3F�U��f�?&<|���7�g��Bx�M��/�KIA~��Ԟϯ�m��츾o��7ze��	���R���̕4���2c��Škg���x5�YTzr{V�-a����W�=tsya����u�����#%KF;�;�W�T��߲�6?�Q�kܝ�3bǄ��JԊ�w�u����vj�f�lfl�k�<�H���o��&�[+^>K�_?�P��^�NPw�iޯ�wݷ�z~!�Ԑa�'t:�%��ݩ�
�D����{�w����w?��x�Y��۷��.���{�������N�~�E^�[�eS�[�����ܖ/����O����ՌN�ы�����R]'�Rf8�~V���:�J���Kb'W��Cv���R�Y>�gq��}[B�(������[����G	w��?���u[\�/FA���_�~Uy9s:����uZ�]X�yoӖ'�����YO ˶-M{�]�N'\:L;,j��9�U4\幚�k[��9	��K6�(ɘ��[���[�bW��K&T̢�
K�={J�ț���:_�lq�����_�$���Z�n�ǚ�U��{G��\��������Q���O�o�Ξ�)]Zwk��:{�݇������C޴�N_��s`��)Ҥ�=�$^��Bz=̱iƲ���<�ƦӯNO�7�������e��= �=��2d�q7f~��HK	3�'��?�U�*ɯ��V>�ָa�R�p!~����3�����ۼ/F��njP#��n/���B������㷔.=�,麳�E`�Z�FcÏɨ�і�
��vtE�~�z\߬�ͣ�������{#�d}#�ʔM.>>�f��ܱ�n_/�D�<|�߽u���o��w�z�<��C �>�\y�����pPI�j�����ܜ���S��H+R�.��1w,�5��z��@]����?�~��a��u��'ޫ�+PGJ�u�٪닗eG����?6�RRެu���&\�~P�������]��ʴ���D���jؚ+�����T��,��b����Ē0�/����f����mrB�����[
��1���[���?ߺzݘ�y��s/U��d�Z�iޚ�q�����Q��P�~�4�F6�]p���F�A�O�KV����̭�i=y�:�������[���<*��J~���l�j�������r�.Á�o�y�}mQ�+%H���>|���⍕�>~��bh����o�D?��af���/8]�vk\�ѩ�#��hRÏ��
��*n�k�3��d���;�e�GO�u˃}u~Ƈ���訓+nx����C��n.��]V|zհ�C�=�c�Xgn/�^U�]Q?uM��w����>1}萠�C�ic�p.tEZ��=��(���*�&�I�87s��!-u-��,���5e�xBz���\�et�а��S�)�D!$��k��j����.��%�/�k~
��ó�h/@n��KL%�Br���Q[>�մ��u���7`����5�M�*�5[6u'�}Y7���珐�ש������}��7{7~���z��Tt������ꠧ�Y[ݿ��1Է���PK*'.D73�	�sG���0�e~�ܬ��w��S��
K�5�ή/���1
��=}��py܌��͏��n�!o�y3�s�2S�����;[��<�CX����ŷel�1��k�>okE	M_q�-��ǛᲦ��3~	�քs��>��H�+�����Н-�w5.)��tt�^�sU�.��E��YtP4ngf٥��f-����Pbٵ�;��9��yw�?�5l��~?~+�_!�*~*\96�ze�AO�і��,��ԧ�;�����Ț�����:���0��`jE�}̩��Ս��+Ʃl�Qz���>��M%*%5��HP�Ӵd���{݉�o-�3p֘�i�է�gOÄ�.{���h��}�;�l��|�z�ݒ�!7�e ��y���G0cɎ���Dj[��vIS��Θ~�Ew$�=+���O]=�����k��V^� �m[����uH�}..|t0��s0l3,]UQ��~� ִ	(�2ҺH����,ߚg������c2<]kl����/���<��8.�x482e�V׎O|eL��t��/���E�ޙ��������se�4�-�]5�Ա>�5�Ϯ"6lw���u��ϵ���R�-+��`V����Ξ�Ztn[��5�m�6�^'Z�xk�͢θ���b�6��ޥ�U)���.�|�����,��u����}�n%�>7��)?�7zR�}'U_�lc3�@��|	3q�Κ���7\���O_�v���]S�_,����)������+2~G�9Z	K_4yy���[��;v7�'�>���v�?��m�/Չ_?}���u���C���:�<1�_�I�d�7N����_\o�
��n;I�1S�ݹ��r�C���t����Y�Aw"DMk��onޔ��k\ű�k^���ʗ5��N�^�Ҿ��f��>kG.h���ưom����\����K���bIל�)�a�3,�1����鑟n�4G�%� Ӎ�7�͆�>C��#�����6�R܉A2{���7=A���������ҟC�W��\Y�Izz���Z�����6�]�}�<N�+���zY�X�Ŋߟ<��gk��X폨} �4��ĸ��N�"�����~R��\������������O�c9{��r��]���T����̃-�������'���Z'*L9�<c.B9\�vK��A I���O�֌�U���%��T�9�$-��Ʈ{ڐ�����/����GV�=�v��O�WzPN�����q���''���F^i�,Bh���<����;��s5c��A�ӵ/�y�t�R�fwȡ��w����)w}��gm�����vٿ?w�N�ű7F���,{6_Ŀb/�##}$~ɸ��UΫ'Vd�Ov	���cF/�t��8����f�ٔ���{T�|O���z�]�V�����K�(^���~K��9t�1��絥�0��;��mY	V��	���N\ޣ��3C$��,*kZ]�cw��:fc|�~�.��[7�A�f�~��~��S���۞GVLSZT�7~��ĵOgwe&�/��� ������7I&�&�[v�-4�In2*��ƭ���0n�	�S���AKƃ�n��Ӷ.{�5�a�U¯5���+K�>8DB��߸���7���6bQ��^����Cߧ�]�zg�M��F`߅�����������������ԏ����ė�3iRIuVn�]��w�~?g���ޢ4��N��cG�g��\��4DChS	���2|$E<N2ka��U@�ȑ{��g��ʠ-[��붏�i��c�&u*�Џ`/1 ����_)æ�c�I�G4��s_E�a/��~��o�-���2�(u��}F�_�5: �U��"�o�_��K,��h=�l�T��I|QqΧi��&\��P�F�}s]U�b�8����[��_x��q�X�|�~��M@��.���.ܞ����x�yx�����8m-?3F������F$��zvq)���b����&m���?�,��soY�SG�~T�#���/����g� c9Ʊ�d~�&�ι���+���ӻ�h[����{n̂�C{�L�-��췫B�dl+Jx�z�� JY{Ę�$���7�Ϥ߹hm*ͱ	�}��l��-?��k�VU.���S3!�y/�<�5N�����x�/����Ǯ:1��YV5p����o'��p\:yg����qO\*��g��G���jZ�`���h�<����ד[��W��&�7�.}K��5oI��;�Wj�\O
���n�	���#�m{�ά�2ީ�����/����-��~����=z���<�i)��UZ��9��[D�c�'Ī�"���Ο7,�K�n��}�/����:1�QFT��T�~�a�eòemCnr����}?�y3��>�W�M��7[�ے�_g�#�~{'j��?<t��H_Q�"x��+�����Gn����|�gw��H�{����������C��s��&�{��A�3�eg��\�t�e���˘�:Ģ��ҩ��/-i��/nFM��zK���}��7��Ö����u���+n�Q��y8�8t(�?��~]�D�����>;�`�5���I1=�ٟF���=�I3ru\��j��%?:q1�_�N��\s(�`e5���"�J�k�,*J]m�V�?���O^������1B�9ٷ �W0&�My)_�L�ui�b��=�O?��� vm�Y?�p=s�;=����!����e-�� �%�"q��a'u_�z��GK?�w@�����_��>6a�!7���9�c�Q�}�����ۏ�^.~�������'?��p..��ϖ���ih���b�>N��S�>a{՝<�i¬9s6+/�(�fv{��X���C�̩m}S��Y�DA�'n�P�0(3my�/@�7?�{k<Mw�Sd��)l����/-zshz"����a�ЂG!"|���U�ۛ_X?ݡ揄޾����-���m�r{\9�=ߖ�oʻCc���&�ۄ}U��a��oo-����ey^��m��=9���ꢪ���?�&���^轜:�F�t��ĉ�%5����_�=�YS`^�k{�R��\x!r)�{f<\�)xh�ǧ%-��O�� EĊ���g&��,��I��q���_�Ή���������|Щo��ۥ�f��jU������`�fW��ݨ�L��\��k�B	S6:
f%L=�U��g�����vx�{t����Vo	�1���nT�����O�	�z���;?�.V�;U�r�BA[e��ϥfw�hr��>p-b��6��S�Y�z�CGm�c�0��+?￾��������"1�7�ʲ-[I��Ծ��9aY��/.M����GC�7�x�m' �?4&Ѷ7�`�FM�В���l��Gq��L�F��|����������=3�V[]��;7���hj�
A���56dו�j�k k|fO*��\�oN����H��x��ͣ��K�t�z��Y{u���3S��5��>�7��v̥'՚]�L�}0�h
�d9fg��}���,7.���1��^���"gS��v�����G^�P7cԝ��a��ѰÐ�M5�ҕJO�=��_)c�^8��Ԏ#��G�\0��C�xoW���-��
D���	;+;�Y<p� �m���h�tlďUG��5ne�o��9�R����4�y��Ǳ��GS��/�~��پu�.Wݕ�f,��3␭KS�;W4�]�`T��>��K��w��'�����7` �۷I�C�e۟ߛ�o��FUKS�tvT�sv�U\e���_��Д2�־j��~o�;�����f�G����H���Q�|84M4�Y-�|�A��N���+"R3�ؙ2�x���,s�z�"�BU%�+.���`��B�5�o�!�/8�=�:cY�1��_��^	�}*bY�[/j�y=��]_Z��Ԫ	k�M�'4��L�?]P�o��-S�>�$��Z�%L�wX_��hrܗ-�/��V���]X|`Pj=�;}�4Y��]�۝XZ��j�)�3�^�Z�es�"n"2��p�eQ���1��⺌�H݌םf��_��;b�ڨ+ш=\�Y�4�h�F�vO��l^���)4�T��^�U	���gG�����۟Ǥ?	�X1o`��Y���Λ��ד2S�Ƅ\+�}���!��x{+��ְ�Z[}��˱���>���~�
�Ym��)���������%������m-U�5�.^w��Ԙ�B���U]��P\�l�����@��S!M�|h,uʓJѾ���/�A��&��.����҂;wzҶh9�x�@t͐q����є]g)p#��GY�㉾��¥����_�6����>og&6m��7	��ڪq��?��#��t��[�[�=B��iI�:�v��,���X�����|������M���ۧ�z$c�#ӝ��)��g�f�N:�)�L��!oBzOX+Ϟ�y�����i#&�v+�pM�ō��|��L�!�7��J={w盇:a�7
��C#�&�۽ag�S�vc(�\>t���y�V}��?L�#.�����x��P��3_8��Ĩ�m�C=��|~�y�|��Uc�j��c�ѷ��ں%sC��>��5�4i���H��~�ɵ�:r�g�2����g&�t�l2�_1��w},��HE��y˫�mgI��S�Փ�\W>�J�	�黧�
�"�~�^�2�`yϭF����chq�JsNo}�<��|��@�৩+.��'�.������K�����o�R��tWn܅S��P5*0���n8zJ?�h��殽���%�;��J,{�����&�D�RgG�/2��=n�@���fU����E�H�K�I#^�pQ.	��']JZ>�0?��ګ,~㌷�Ԉǘ��o�^|i���Άc�a3�Sf��^yC=i:j��_�7|�n��:�04%<u뀀��v9)?�-�����\�8�>�@Xpa����QŗKW0�֯~y��C*�@r%i�'4��y�=3e�-򐓆�}>�C�E?\	���Bу������^��{r���T�+]�uw�����M��]6��bG?Oŗ6�@�I�%��`<Ո�tp����n���v��cF���rd5�ݬJ'L-��X�H������U��9�z�b^c]��'�g]p#�zϜX�$,��>�R���]j� �vkHa�r�]�KJ��P����i�����邞�������\e�-��d��6D��*���?���;���(�o���K}��͹�0�zl�8m�c0õX��]�f]M媈"��t3��N�Ӹ�a�U�OQ'��������,p��N�^L�<���1�ۊڐ�����)]{���y���7�"s����cW�iE�E���`��P뷤��O=e��Nn}g������,���ӣV��1?�`�4ce⮙cGx����ZW�����۞>YX���c�ĞK�NZ��t�ӻ�/�-{r���EWǈ���'��9K�G �&-8W�K�=���]ʠn�����o'/>��3���E�(�W�¢[���~�����^N�u���E���O�W5�>Y�]�}�w�u��D�����C��\!m���r��?m|å������������e��<CH����BW�xߐ㕙��O����S�����u-҅����]5�8Q�~<�怤�U8r��������U���=�_O��Aj~=��es��j��������^�YYHz9�4q���]��/��0|IHZ=��mJ٫��O�S�{f��r�Ϙ��|A�WF��4[K��<O�����<:J3�v63������/��G�G�]��ga�zs�E|S�zu ��-�q�5Q���W���.�~<{q�OE�t��Ʀmٺ��@)ȩ�L�#�(���l�"AvA�.&�H�b����>B�[�w��/lߐw�դ�;��+���2e�U��:����H3�;3bF����1�1`y]�xw�s��
p%���Ǧ�A����W�'����Xѿ����q����F~Ǟ��5W��x���d��^7Z�����/]����\fm�[o�E@��I�HYRX�D���b�z�CB\��V}��i�>��Qe]#:�_���U9�jqҮ�q5��㶧]����f���Q�H-�T����{d�A�L���B텢WW�)o{^�P3��[Iq5�\��Ts��т�٫���'�|��,p���R��w���C�=ҿ�w<,��;cݨ�};���Y�/����6��zӵ�_Vn*�=ܶi�m���+��xl�/T�r�֜�1yK�T�[qb�"i^ߤÉ�_�����<p������@V��X㘧�w�A�O����I�.�����{-P2�W7ld)t�i���kȭ1y��r�D��R�:f순:��9=�M�{-ͽƌ�C��8�k���Z�=�-��Lr�����GެX3hHX�pЌ������.����!kވݹ\0t7�b4�lGx���sO�f�z	zl��z4��4����ç#$����H�b�/��<�=6����k��=ِvi���k��\�Y5�ք�Ǎa������[:H��	߽�9�q���	�a���3y{ȷ}��N�hOk7y�s|�@V��m�������h&v�6w6�:=j̩���4��G/v͜��qͮh~�y��jX-��h�������\Җ�q���_�{D\lpFi	�(���Rpv�re��	b�����߹r���[�5���s��x��+��l�.
UF"����7+���#k*��>��Hw�p"��wc��_���ִ$ p��E�+뻴-�æ�[�R��<��:eg�A�I5��߯��ܮ>Io�U�B>:o���2?�ە���5�Q�ls��pcW�&��޸8f�s�г	'������4o��Y�K��f�d�BG�6vz�za㢸v�9���e�!��=��B�%M�.��ѿ�^�hzO�Һ�$��ǃ�D����(b��*Muq��kYe:�M�!ν;6z�%
�׮�z~�ʅ����E�Q�{t1k����țD�R�j��.5̥*H�=g�ʺa����s�_wo-����Y
�l������uߩ���'%�i'Z2���������L�s��hߏ�I�q�]��v�Ɠ��f^�8H��yp�m��iC�3IȂ����g���<�|����C/�z���%�2/^k�@�P�C�)(^�����f(�d�m���ٿfC��"��dB!J%��G~]}����M ��eSKȊ2����M���UK��A�8���:�P���վ�nCm������]���d��4����a�"5o��|�{r꓏�LE�m��S羻�j��!��'n�-��m(�xz^��>���BJ���3Ei�}�W��ε1���u;����ʊ�V�/y�u֯7G��6]��oZ|I��s�P�z��ʖ�Q��Ó�~|��=;�9�i�+�L�fܾ����ػ��w��g>���/N�~q�~Ƞ��E�oO����Xw���E��.{�A�O�Z;���C����p]�h/�%4�Ǒo�{�(�~�H�_�/A���AtRnq�ܺLZ6��[�~��ҳ'�]����3�n��״�q�N~\ԹG��#���2��A��H	�O�/
�y.����@1�ޑK��rʔ2��?2��G�?�J�3G��+9�SF���ÊSiud�]��3�
�A�V�����w����hv��F���Q���s����s"D�`��,vUl:d:d������ӡp0
��P@�L�f��3��%!�ȳ�O���E�i�N� ���L�@�[� �FA�?b%�9|f��;���w������ovo���rF����\�)�n�����T UF��OJ; x:��3�G)3��I挑Y�F�B�����pv����kN������{kvL��$��+�z
�*�(&��^Qԙ4�u��z3p-rZ�|��ӱ���P�?GCp��W_��b��>������i �4�P x�1��O���\��`X�:������T����4�I��e����e��e:����w)1��k���7Y��Y��ҩ����I�����JZ՟WVǀ�����t�����R�������?�����D�0��3H�\��0<�����H�! i�J�/#�=<���``����0?XL�������p�T|8, ��D�B5bH��
j�C	��pX�����X����H�8����h�x����Xh������106�b�>���9��P��(����Q0��$Ђ��p�\��s����_~���@9�"0\����2���p�����ѓ1F�!`���!b<R`Z�8�!0��9����3�\`��yQPp=ph ��pp�c�	23����H�R�!�D�t
	A����X���ѱ�
�d-�+աp\��M0r�\��F�I�lS�1,?S�H�|<�E�P-*N��j�����@B'SH��}0 ��W ��I�"�Q&{�b#Z$�h�2��!��(�4+a*��&�j(�����:������z g��F�Jb��h����N�[i"����l.�]�p[������r�p����3-��x�(�2��ԫ�|Z�d�A��xLQH�)�?��k�2��'�I�t��1UT�ƫ<��C��D�NiPP�����4ֿA �_K��� �����*�*1�k�����j���.9��n��F�Hd��&�Ka�"��`���6��fC��v���G#T� 0�(����_�~i�|��I!�Il�ݦ�J�2�YGR�Lv�Jg�9�J �I3ˉ��X�
0�k�dr��	4�к��_�h=��bI�	�Z8��+dA����Ђ h�[΢!�B�f�Ap�"%Yx,�g��\4��(��V+��W����6���D9�F2b�B!�x� ����N2PmU"�9�AY E�癑&��z"�Bo�wY��
!4����3� �a��vL�aRL�M�RIj�Z�v��F�T�w��d �@�LW�q�[ !B�R��	V��n�Z�������t����'3E.�R�y�9���^/S��+�(cuN� �q�l��ĩD>�����t�ZhқD��oE#�*:�	�A�)�� ��Hǣ���u6������7��i7�X8#C8�\6��؁��� �u �ˇȴ^!M���E��"���2�n:��Y"��cs:�L���#80�4T�Gc�۬`�҄6K���*�
�p��qu(}��21b�����2�aW#�T9�G�K N'�N��2*]k5�(����ىh���I��Ie�Y%~���5�y��-�J�Q��Qt ��F�!�V��*v��������wX�"�U��ۈ"����A\"Q$�C�\�!��h��+��P�� Re>1^�T�p*J`Ax���`�7`|^�M���|�S�bv��T/�H�V)K�U� f����P��M�(]��F���4��(���@i2���Mp��tJyz.PD�v��K#rp6�Qʑ(���r�0L6���|�OƗ�1.�܅t"U~��3�H4��@YB�R�E ����Xe�B�����OŃ����3���8[��Hy$�؆EX���W��q:\fȃ�� f#W��r�R�_j
�@���c ~:�tB<6��f�y>�)��Mz�IVp58�����ȱ�,�#�4�F��<`���)�E�q�<L��u,�s�o 2+g�p�T�.�<�<�ΎU3�p�hG�(	������<�̠��*����ZKO@Jl::^�U l ����RN8�`��Z� �(�R�G����beZ�)�Yy+b�+ez,U��(��]��(N3��)�T��#�9D��a��_��R�*Z�G,����y�j�2I.���CeZ�^g�1ƀ�K5:CFc�� L���v�k%z�$���dp�n��eXY0�N��q\,�	|��Ʌ���nTAY�j�� K�(��N9�(�(�L�t.��!���C)�+\�P���G!�2�R&�5�Up�A��X8�M`��6����`��#�p�����B5�� ��<�'f:�^����J����9`'����:b���$:�T0� ��0��MdɅr��
8&(�a ��;�(�����
�����,�t����.��f��P`�TctK<&���p��Fa��$
����l(�#V��B�Q��(<\�$9�B˥�uL/�9H�>�g1Pen.V��p�Z]�e���RΑ��81�Ƒ�� ����(t�����3S� ��VE���~�/�� h+I�l��#��u;��`�Ԇ�p�Ȑ�}H��.V:�*�Ճ�|	R�B0p"���@�j�kI21�g�(�����uj#	
���N$	� 2\v�sY=P�a��lb�	*�)�>-����,� � �� 18��ѩ@�@Bp��~,���C��D��Er��dD2���b�/gQ��Ah�t�3)x�O�Df�@�|���m�_*��<V����0�L�Sa�q=F�MdbX�r�,5ҥ������)�^y�Kq}>���y,~��hx0+��$� )�JLB��j�Q}N8�B����0�����]X.U�Pf�Q�B�[�S��
�����!FY�r �M�����T�+d8:lY���b5@���&�g�u6�ͤG��E��"%�Mc�,J���rl���N�X�v�ɩ�Y-[k2�|T�L-��l:�Q(�hHJ�+96?�$�ZF��� �XH"$r<X2f�W��Dc�D�Є���8\�B�E��6�L�{m<�ĆB�P�M�"�1������v�(��d��`P�IN"K"����@�� `�p
<9��%��1lN����L����B�P(ū(�	�p,�Η�m�
�h=��J�33�
�WFH��Y�)(T�' E"�]ś�n��y� #U�X}D1A�'q�XP���b�H�x0��I3�l������!��>���R�0�$�xY�^!��Pt(w`��~'��H�+V�:�2*�i����FD�M "G�0X��qEN��&�i=���I�>�B���U�@�nˁ����ݬ ڱ(7�LU�B��l�	0�G�	.l
�� ���&�W����D9�ʤ��`�_����FG���=��(��� -�-�����0�6�U����J��!F�8?���R(v�ѣ��Iz��*�q�\���r�1�w�
��@�C�4�� h\ 1�>�M@�('	dtѝ�Q'��v��@wX���h��B#ج0���W������\�6�x �Pbk�2&UJ���$ ��rLN��`�8 =� I�&�q�e1��F'J��:���l�1�$KD�؈T�Ǧ�!z�=��W��C-hl�g
+� 	4J��eB�&,��0���v�C��*9���1�\R�
5@�H�E��V#Gn�R�*p (��h!*�]tB璈�6&Q�.�$3�j�����l��wf	t˄w |'Xg��IH�rf"@�&�Ni�a�T�R��r!jQ%F����JA�/t�[] �[\T��
��v#�AnG�JlP��N�Hl>�	�0,@�Ƞ������"���~8Y�t
��TKA)t>�`��`9ՋP8$$�Rϥ�5H�Oс�P$�I� �@$��~9Q/cu`4M�s�0�Gňj���tl&C��t2�����p�T��92JD�,A��:
 Y�8���p�'����� �G�T�d1��Si(��kT�t7	�pqX�]�Z8-C��:e(�W��Y��"R	u0T���c@�N'��B�J� ��lh���$
q@���V��h��|�k�Hɜ�W�x�tg�ot�%�������.S���w"��':���43L�e��:�\����
��@{���%:��C �@�N��!���
O��M�C�%N�� ���5	�<	GG�����8���Qv���f��sh��4x=�$��i����d�ډ��4��� SΓc�.2*Ј���X�:>�@�S�@�K�DP���C ���B d�bC:-H���|V�U���N5�Ȗj�X2�T/a��H\0VEuٜP���F	����W ����^	p�b����8�")���t��B7R�N7_�WEJH�`��.����|��&xu���4"���T��t/���������t����z4e��2'�����b��YI�x�d�^ �B��9 5l�η"��KW���\
���L�V`hj���� :`�b�ڀF@�z��i��UVQ 	2��q́���vL@�Yj�`���c��}���V�e�Sd ��~#�B�
&,M'�X�:4WE�r�x"�
����� ��1��T�����"
@9��N�P�l�L`�4t����d��@>��`W��u2�@BA���C��2qb�N'�t��e�ڠL�&8�Xm@�P;A\�TIc�f�]γ��J*��6H5�ŷ��>	�#�L:;�)B�(�̈%h�L���0����R�sX�� eR�.�!!X�p1������;�D���z���(/��[^]�ay�$ͪ��A:�� �n$@tK�v!OU�I��"0p�#S��,RbQia�M"^&	�r��
u���+�|� ��!Q*c`хt�Xd�PnOܡ�VQK$�9>*�Uq��W��$47k��v��e"=���e�df��	�y
�W��UJ6D�&��j��@��*�¥J�O!���-�=.�DDO�����*���� L�Q ���:Mˤ��r�K�1��|���p�
�Ii ��<�:��hy>�Tf�"U`� ���R�n7k�X�Ѓ1D�f�B">`z"%T5ډ�j�T��F���2�0��@�b�$���b�\�PyD�HX�@d�I0���"��M�KI.��Õ�;���hK����b�0�X(U�s��d���r�H���W�nu �B�l�S�a������$����_�&�Q�$Z�z9�J�I�"��j�E�^�$��v�\�vpB���2n��13`z�a�Zex�@�Ao�<�HC'�nMl2���? �g� :1췺�8V�.z �px"Ũ��4�+�:!E��D b�*SH.9_HG� (��]��+�\8��\:��Cj�R�b��$`�õ�`��aq��!vxl�Ds�P(5
C���@Әh8?�H���Ǩ'��*HD4h�z:�&�Ӏv��aA�$;* �|D�@���eJE�]I*��b '�C(4iLF���x�V������(�!� )Ɍ���.	\���m.��"wu 7�G�1�t��,p����a<"O �`�B1�#�	l����k]���Щ4�S%���6����D(���qe	%�C�:.��1Y���)��g�i8��L�0,�O�@�L��f�p�"AA�i)#�kai�\�(t��
�/M�s݁9$�������f���䁝��Q�	(��$)�TJ#�S�65���i�8;M��!�d9�J�Fˌ*�F �^/�'�Z����������(@��t�gl6��ƊĀ��Z��%�����<2�4P����.���|�R5�T@8`����A�P?�!�F��zDHi�s�>��k�C�j0��W��M�r�8M`�B4�٨�D#@�2�@L/��`}1��0l"��LFqB*��CзLEJ�pنPw\f	P=!�6�qZ�Fo@�h4n ��0�%�cl��z�K���JȄ˝@�E�+i$��cAv$h��Oe��D�L�Xy�M� H������'�I��\:�Jg��8&"�1�zJ4��ē�顀 �"��B�E\����p	�	)�1$������g�B��2ɜr2�*��3I-���<���O\VB8C�h<��y���4������yh�ˮ�}>���sX�:� +��4�,��P,��J�pX��!I���s�@/��3�H�͗J4��t�3���?J����D��&Q�:G0s;Xw��2v�/���Gx1?ġ�8F��H���Q �eB��.�1C8F;^�`�� �shD�W ��
�`�h�AǓ�F$�s�"�fG��*3U�4Ҁ�P�5�گXb�i�
p��Ǳ�Z׬Tk!]��}al:�[�����`�ڸ�J̡�0x2A�l`���a�~�H��E�q�4� h.�EbP:�xm��#mf��k���N�	
�� ��y"����	�F
�
d���@;L�Yg��dV.��ƈ� =֤�Xe/�� �D7ʬ��l.�L�5��x��p!i~J%��h�����Lբ��-:Uǥ|�	�31�Nt,�Sb�	N������ ��5�l�Ia�{l
!� 1��r+����iV;��0�}r0F
3�2P3{��)>�� )�J>����H$��+d��d���G�t<�P���l��H��lNs ��4�ڍdy5h�(���,����3 >�M�4I�X����Z3X�6������]C�1,0*���>���h�.����F�r3�t>����r�6��&ErY�r�X�@J�X����Pq(oC*46�(��J�U���C�!\̎9������zER���� ��k"��N�g㉁f����$�� ���h��HUr]� N� 9�Đ���,�	Њ�0�X��c���'�B7 �yr'��@�}8��(s���1�:��/�DZ'Z�%P$�Ƅ����M���:�[�d?��z!L<�
��$D:�!p�/w��l:���]=��01�	��I0�Nc4j��"6J ��c"�4�g�Y]D� �L���2�E�u�\ SY� �ƌ'1UL��$�IT�W��;�g�`�DC;B	��Pn&���(�UαRmD��3t<��!��d"\��8f1�3ѬN��-���`��Bs`F��/�k�6�L���ي�1��|��Fs!}`,�mB
�zK2(�\�IC*̒@���\ ���{=<���F�x"���B*؁8-E0a�M��P?	��Q�@B.�)�x,��v�7 ��M-(��"�@j����X
��s� �L+�bh:�N&0x̨w�)x���i"�$5w�l�;-$�@*��D/�d�~�UJ�ʸP:D��E�c�(B����� ?��TV��-^<-eY�\�L�1d^d�`#B�c��|��Ŕ��`��E����P��,��S#�"�����F8��
4@������_���}��t�����"���22�j�HC�}ZS �y�x�P�Fy(��KU�?�`P9�r�����F���40�N)�j��Z�d�84��W����[�hخ@PU8�;`g7�@� �R�g3]P��*F�=.�d�ٜv�I-DS��7�F&6�c 3�,�i�r '��n�Wh�lb"����׹�v�w
�B�����KJ���X,S�` �Y0B!Ƃ	�t��7dqr��#�H�\�#�b��8�(�	�� H�(;�..��xB�W��t2O�Ã-p�� t�
Be�H|�@MDw X!Kd�|6�Ӯ�8%H���u* !L'�L2�I2����<��v�,@��Ʋ� L���tOO�ZV�ϯP�j�d��}
&؂��a:Z�� N��qZ', �9^�+$sh6�v���+C���W0�d�1����*IDG���!^�`�$���+\��������a�p�Ng��5x����
� �F���n%�H2dH���	���
yl3�#p�D(�lu�P��{R�8ö�<zQ����\��-Ё��  	t7A�cC�00�NJ�T��3�6�n�#�D�g��X�s0:�($`��2�B�W�sW�����(���3Y "��trqt����R�� H�EȂ��N�����;�	���F_l��&�Cs�r�ш��05O��Sh|*��������@�|�S�`�G��9~�W��C(D|@6�h�Z���b�m1iNG���cƈ�|5�XN��iy�R���7�X�������᠁V��Ft�ehOE00�
�����6;��;�xE �J�J� ���ȀOg��$�����"��G��%� L2HY|�M��r�"�@,��-��Ut�	E��Z��쵣�J�C���(�dt�"ԁ�'��C�`������m#e��f��U\%n�u�P��|/G*�q���h\A�S�Z.�Mr�Z�Pȱih6�&@�1^�����@��?��ԙ�?VBT��C �CK�]<���{*�JEe���m6���f��P8Z3�e6ms˥X�*t*'�H$	u�K��rO)R��:��n8�W�s��8�������wy���}~����=^~)�
V���A�jC+^{�g���������nn�VAs�����%9����\COps�^�%@�U ����jAӘ���>��[���:b��5)T�ϩ,�'��N���G�P� .��`il�d��w�5�œ�����b�>��T~�Ƈ�}C�P<�a�t&�KaR�*���/�PW׀!a(�a����>^_OC�0����':�~/�9�����������Y	�E�zQ؀�3�DG:�0��*�.�3��U��#����C5p�H��kfj�A�1:S=ԁV�m�{#5�E������W�z���&d
���-���H����סq�`K�����p���:�k5;��ϚYl�3�Ia����ր#�H�6���zx=��Akh��>���F?�u������A�dM��	0��������5��09`w8#�Mx�We`x����ї��γ�qkS8���#� � w60�l@0#1��ƚMar�e0�>X<��N� ���̉`����~��%�$P��MV���ׯgp24��hU$����C���7��eXF&��5aR] N��4h���0C�O�p��)���
�M��1s.�1���`��R����G׀���>�u��m��*�lX@]�?P,��_R@YD0ZqA;c�P�Ԣ��6��\T`�K�}�L���������K���ׂ��#�E�_�m��������!B��Cy "�"z����hp��BD�+0���Gp�>�Bu���rD�}���p�.Fl���7��ۏk:����h�c"����~L����_hD<
XX�7r9ñ�6����Np����p��H�u@�G��/+sc9X��i�����b�ހ%ZZZY�JrG�� I����A���ڟ�_�[
��2T����*| ��5TC/��
�Kh�|y�yi;G�82Ƒ1��qd�#��m(� ~����6t�@�����>P�%H������blD
`W�K��+��6�� �nA�o"_��X��nX�ۣ 4�c��@�D�����180=q㿅L�8�cc`��o�R���-�P��/�X�;�?d_�c�@�"�7�7,����������6u����͸P��T���@���;���8�[���@�1���NƟM����c|'.�s�Qa���Ƌ1�
����-�A��@n`��hb��n�����{��8<V��{Ψn�Ӯq#�Fƍ�72nd��?�H�w�L'm9/9�a�����><���jx~�?��I&Hbs�8��w�A1j���7�Y8n��}~o�K�߭܍a��l�UUx��A{��6݃��[�j������
���󽭄���t��]��sxj�^~�ڪ�e��D+�Y�L1X��~*$1rzMʝ�G�;vo<s��i��w-�\�Au��'�������Z�ݑ��7�vl�%W�"w�k��}��aVb�A����K����P�!E��o�'����#ME\J>s�����������#��
M���u��g��1�,.�^çY��XL.�|����Y��,o{$��C�H4�JR�����P�K��0p���t6��=pp@K���
�Q�c� 0X���7�ȊN�b��aH��������(���P�����A�լa�uX���sc�o��~��1�J�l�
�ګqx5k��K��6�.�7� 
Q��*�~G�H���,~�!�0��a��݌��p��QP�g�����Xu]"�9����u�����p�sH�TG��$��g����W��]y�z����v�֝r�*�x%����c�I���o-�N�|�9m��x$��&m��-�n����ɓ�_~y&[��}���.��e����J���->*�Ǌ��I��Px��ēO��s�a����,RD���&���D�G�>��.zuN�VQ���[��W�k�J!{��v�H\�׽��M����-���Fp�|9m�_��3ӄ~�|E��m�P�����Qi�D/�p!����E�{�����?���R�'O�b��?,��4����h򦞪��w��\���Fv0���zm�������ٖ�3s���'�n�$�I���%�%K��I�E�6��]����c�=G�����1E4Q,�J�QN���R�S��վ�%l����e�ֻˍ�e��ˌv�������	����"{����&��h\{���Z�����Zr\>Y�X�_TZ�Quź.>��Tmje%t�a�e��j7'D�|�)��:9Tu�E�X�P��t�����8�=Y�HZS�a�D�b����kds&�0��R��e���7�Yk,O���ܲޤŝ�nwzj�z�J��*c*���2Z��L�%[v,	Փm���PG�(�Ahτ�QIU�B;"]�^�����vY�Jc��C��	q�!�2&�uB�x9�(�١a,v�m;�SW�X,>�;mV zm}�e��5?A��q!k7X�6���M���H�y9Z����V�T��x����|�a��q�rvR�����]6��J�A皺�J5��w�=�(�ᆿ[BQ�T�݂I!�~	<o)�h�ޒ���L�P?wbD`DGu|I�������ih���īM�3�?��՚�+�Mv�9{G��.lj-o���ƽ��"����0'\R�������,�+~�8#���nE��M[�x5��T�k�&�$�'�N��BN⭔	������S�?I��Q���Ke�;�gN�������J1�;��h΄k�E�K�.����!�3�ׁc�WF�l����ʭ�n�=�7F���]	��������'s31��S������?�x�R.��"y�뛮Wl�,�P,Ӗ��╍"Ļ�&�ΐ��Mt��+|b���)Q&�,�*&o���mk ֘�F�N����>94�0��٤�*��RvM�m�ڽ&i�������Z��D_����3
�?w%ejޮn�K/�-H�m4�rNM?���]Ȩ�<��{�ۏ-�����G�}kS3O?����k�&�P�{-�3�o$����n�2��:�Y_��5Q���{���G�w'y$��������[h��=�>���m���&j�D�{W/Z\���k��U�T|���ob��+�f����d��8hJK�nD'��I.R��[�`��k��BBm��Fٲ0:Ҩ��6�CX{�����1��O����p��<z�ni_G�Ĳ(��<����r�awH��㦗�aE�ֻĴ#b?�Q�����D�d/����ۗK���OM�C�p����D�`3�8�hE�f�6XIF�QF�l����]	ydq�l%����W�ҏ�/�H�׽&p����z*"�r�D�"K�B�;R�bN�7_|���tJE��4�I�m+,�	�X��3w�Ve�j^r�����x�%���M�<:���}ݎ�6U�������͵�6g�L5��<;e9����e����L�0WX����r�m���S�<V0E$"��jm�3�گ��d����V�[�j�R2
^{lzSD�~W�=8ߢ<�[�h��!^<Ҭ��_VM��&�\���#3i9pNI3k�5�C�$��6_�r�6��MV��7+H�N�E���,K�ڧ�d��5���O@QfѾ�V�����u�kYV��x���5��AH�[��l�I:{��%ᡕWTړ������0���_U�K(ǜ���N2��C��uz''��S�K�>vYhU�}zH�_�.�A�;�������ۺ�IӺ%�3q*�>�Th��_�.,��V�(��0�-���:����T�\�D��;�����?z�*ȿ
�{��@h��u����d�u�Ԯ+�t��
!<7<W���:�'w���,�4�c�?����!o��g_]���A�C3�μ�?AK{�ْ�ڄ��_o�w:W/���*u��K�'�Tl�-Ͻ�]��!��h�(��|�:߽>qKR�ZS<����8-���'�yȬS�.�G|O*?��BC��_�S��ڶ�G%CB��_Q"{�*����V9�(����L�q�;Wd��YzTDOT�'h�f;%=-fe�x�^ø>��\�L?!����iʤ���Br&R]�́�ͨ&g���]�n!ef�J��i�syx>�!�#���
s�Ċ�*7q���/��s�����}���klu��d.~�$�d?�&�ǝ�ɮ��\�Nl2����Q�o�2k �}i�wS;�w�������=�'�m��XӠ$�K;��W�����7ɲ�-�x��/.å�m��-V�,V�7K��H�����$0wZt[��ɽM��=nZ�����2�U�a�ּW]/�|h��{-�kI�j1�����_S�������&M��	$��$MS�_	��%g]~.p/ֽ��9������29�m�][NٔFȔH\j^�a��C�ʹ��&��`<*����ab���"Ü����J�qr9���%�4Z�<\.������iNju�ꛪ���7�6%JԈ}h.t]��[�xbK�X�=G�U���V��=�dfV)\J�/+:F�.�V�I���T��7h�=*c��к����G?�Ԯ�[E.z5�ܻǖW%r��qծ5~$�Z�1Y��U�M~-����W3��j��kE��1�fn/mR�R�Zr���0����ӧ_y/��>T���������O����������mC�������R���+F���)xRñ9�ߟ�L+�����/��S��/x�����~��g_��5����ϻ��W�<���m�� ��2lA/����m�>�53���2�;��q#��� �x�h������Z��郉'r{��mfp?b���
�#�� ��7 ��Ķ�?���q-��<�(����~����c�����Ek����r34��w��'mW���BjwE��p|�[\�2�k� 3waZ@��s�J�!
{��+_�zy�ڤF��w�ܽ\͖ҽÐ>>a���*(uE:W�^&�0Ѣkڗ����⚸��V
s��9
^LOe�-�!~��R�I�o���!s�b4�ʊX-"�֝Gۯ@�'H>����D��=fl��k�w�n��rD�<0���W�T���)ૡ �����Ox�V<W�x\NX�k)���F�4.�'|�gxtӪ�*���4�A��B��w�~�ߏ���ˇ�܂�[����u�[�k?/a�~�ۿ����˻�������e��뚱琫)	j�A)k�����_�}:{����o4s!(R�B�U�5WAV�d?_�.��=����s�@��|W�{yU'�9(X�s�����?s�-)�!����/�">�=䥴�PN�T�D��
�$Z�:X7h���c�'<�lL��]���	\p"ռ���ϗ᱌��6u��E�˔�=���G3�U�,q�0}�o��h�L����.�T+�9[����<��C˻mW��H�K���ʤZ���@�X#8�ǡ(�MDv��E�C�� o�y�)��dE��+"ɽ}Ŝkά��zv{+�ő��VFC�<�a7Y(��p܉��M�;��H�������Ԏ@P¸�S�����N���ƆE�z��qm�5�$�r��9��>G���ɲ�"G�nIʖ�+TPk"�����)@��
�ɶ��P�r<O����;}A~������"�̳!��⠅��I
�ttG�&��!�+��W��̈́�2��l�t~g��h=d�:b/����.@� 1~����
��Hރ\��臙%�Q�Gl�B��r-�vfC.'Yŗ�A�;B��lM@�\=0h��{AZT�C�n�O�:�o	c0�����3Ģ���v�K6B�� m���K��-:�W�-�Ɠ=$3L�4c��	�3��'(��ƛ���[*�����E(�$��AT�-3�Al������V�L}���Q�V&0y����W��=rYg澜���A�^�Ƽo u�a�~:J�� df6N!����������Q=�4�#��	NN܉�:B!��	��2+f&��\�Uŏ��^���▰�0��ΞP0��L�W`#�� �{#�	kg;�3�:�L�RNm/��匀�18m�� ��;��P�U(#闁�X5���p:��UZ;Uc��bą.����"��;_y�g?�9O��%��Nf���Qs�\㧍��K�ĥ�#��]���R۱�����H_qݼ��@[|OSI.,�k�m��Ik��"ܝ��m���Q�wҘ�,<7�P.*H�N�Lڅ���k�A��F�g�޴�P8�yӷ8���J����C3�MeXÜe���M���=�̵8I&R$���"��$�L���'�=R?���!���6�Hui��c	}��Ǭ��Z_�JeD��՞���PHMT,��m#�t�k M���:�U�vm/g��~�&*si���������済�N��U�C�%�v�pl�MnԖ�q�ʗ��x<&�e&��г�Y� ���ڡ8;D�5Ֆe�!�Ѿ�8K ��A\Bz,Sg�u�aݵV��=-�C��~��xc�|Ƿ-�jډl$�9`H'�B [w�C��ܸV�m�zh��C�1蜍V��6��b����t�﷡�T�{`�f���w�}�1��)\,K:��@RG%�PΖ�,�xe1��J�5��� ���`�+�u����:���ޞ�_��I���a��U�g�S��"pzl�4�<�7��|C��4ĸ�K`iRvK�(��������q� |*b$n�i���{�#��d2�QS��X�J�G�A�қ�\����(�q%�s#�VA$rF&":6X�m
��c*l�`�����c�sb?�U��$�Q7�*`�\�S=x�e"Xi�X
3�o���p\bؑ��^U��I��$a/4Z�F��&3EF�Fd �"����1ס�ē�Z8���#�����ش��G�<_��]w�o����s���Z�2%K����}FU����4����yg"�6�/c�cȁX2��Â�g��6t4pd$����2���8��ZӬ�sWߎ#���.	���1�܄;�05�=�8��Ӎ�P6FXL�8�Iq��b�c��� �kl��M�ڱ�~��N6՗��J&[�΁�n�!P"��v7��Ü48�Щ^�Lr��ҧ��[�6A�,(�9j�3F�GC(*���0Gp7�#ݛ��+v��EO��{���$�������S)�i��1��a=1wS����ZϷN�A��5Ui7�|��h�Zc��w����q[ǔQ��̓�q��6*�(B�� ȉ8[�z*�c\�e-��|���^C_�J�:��NU�����cK�����^-�����x:c��J!�We��B9�@����e���JBYIV9�3��O{�d�u��}N�H� 8�'����@��Z��l��O�`CU�g2��v݈�����ѡ�.���ɐ���[?kg�9��6au�����Ε�W��D_^�2��ǈ���L�m5�pM4�q���<����q��)M��ZE3�ÿ�S�Z���"zlr�i��'I�|�����4���P_�t��ٞR�$`���]�����u��l0k���gd7�ՕH��6��&�3��D�ӆ�铢��Dv��?�c���n,�-���lsz�o���`�t�}i����K���� ��+�~}UH�����Ǌq��Fk,O_���NO��Đ���S�6�F}�WzE���Y�����x�-�!ީ�[b����
D�O"�>C�V6$M�y_��C�H� �j����K�y������KM�2s8��riYv�l3dS�I	����@����@6mSP�vj݅�yV۩��
j(��> K�`�3X�	�����CC{�,�kb�9E����.Ӭ�9��'ͱ���8���'SZ�7:� �<g[�sٞpiwU�#[W�}c�1ŏ�Zq�S9e/�^M�I�������<�c�j�$�g��6���c�s:��h�%�+�y`͑�!������xY֓��<R��s�hS��Uz~_���j���T5�)O	*[z|��Ţ��i}RK�˧��� YZ!?�r?uk�1:G��9҆�F��Ukc�:x��Ns��5�Tݡ_��s�
���є���<\+���~J<?�}>��X�E��������c��s��Oyo�y�����O�?��^t��A륨�|�1�i�*�hpw���Nf2��:?T?��Y�|���X��Of��]�:�p�8|��˝��鼇��
���٪�����#����+�Q[��k����QW���-��yx��Y��s�{�T-՝�PNۇ�`���er�dL��>\nPq5�}�QN쎡�o@`z����&��7^�U�U������E7B=����)uM4h��\�u���oz����֫M����qh?��6Q�Us*E�G�Eb/�c��s�Nyy��`�m���F�0ݱ+��t�}�^��\���~	Xdh�|R���͋���yѴ�c��s�N��\T]�ؙ��R����-3�2�c4�8��x�j�$_��W@��i��!e z�4
��ζU���u�x:y��
-5l�$��H����#�+�����ũﺗFj!��͘%��/g0<�봞A���L����I��\/�#�G�i��u�~ia�e7�7xCyY�T�[[�I���Nը6J�m�f��W���-=.� ���C�v�����=s^�W,ƽñt=��������a�����n��r+�yw��1/R��i
�48��{�B]f3�ɚ�<�ڄ���/[/�o覵&d,��,��R6��q,��<B�L����Pܒ�(�_��X�XK�p���*� z�T 3�	���� X�$��4OYf<1��Җ#�2=A�d��#��H�Dc= ��P�3�S��L��2�uW����ۺ�-��ǲ�\�BM!i�����%j�ЉQ���f�����2��	��;X�������&AXT�U�8x /;h�=��9�{P��㞣�h�$�$��Ul��t���dc�m���6����j�u]$j���jn,�qia�0T}�5"�C�}u3\�R�?��c�|wM��w0�}ã�uaٖg�T=�_j���yڭ�vx|�Aw r�y��W��	l���;	+'f-&��1��$Ph��U�˄�Q��os���k�W��I���~�=q���g�j\��N]]��T�� M^C{F&�!_R�N�����޻�\9��_&��❣M��f�G3�q��+֐~Z��,��B�(��g�����댿*�&�V�瀢���M��z|�à��{*�:�璌���x2&L2��xSc:�V�m����
	|5�U�á�.:c��ogIkS)�
��{
e:P�L��uZ\��"�#�r�H�ӈ,�g�����>J����yB}A|J
mh{gfNG�M<�H��n	1���rq�z��wfD��{<����r� �6�5���[+��e�l�s��
���;ߏ��&�x��[Q��2�x�ທ���6V�EQ�?Vץ�.��>�qt�l݁� 6��&�~j��(p%Ý7�ߌ���<f���Oj32Vx2A���B�z'[��3|/�Q�O��:�)gX���"���r���#+C/�)|A�f.{/^�")ou�Ȕh��r�����xMIF2��*X�x�i	�P8���f�F��`Y��~XK���Z0A)�;{ �_bgQ|�%Ԥ�����aI��&��Tz^����1ܳ̅�����Fx�e�p���� �Fs��q��N-����A��L�g�g^�Ѱ�"�4�!� ���u��0q��1|�)�_�R�.��>�>X̈,������f
p�v��)�1޼5����d �pW
߁�{O�WȒ(�h=v;��G��I�V��$����>#���rg��QDQGB&oڧ��S��4���$�U�F5����I��J�b� ��3� t�)��:��vulW�k�Y�w�g��>.�����1^_����#!���=I�(0j���4�4P�\�.ദ��%�F�X���@��WjHX�V��^�J����%NՀ�ez���vY	,��3���ťN���#�kw\�#��J{���pJZv:�k�k����zZ���O�n0k��vU�/�\�'�ԗcl��I�x?��k���ۢ�v"+/Ӊ
��J�'(a'?�R?�rjf�elq��h ��Eǥ��A-كŗ�`s�n�f?����V�^V��o
I}���|�o,�+z�/ފ?���i�}���C���ک�;��%���ɍ��P����v:w&4�\
�&��W���z)8���~�-��l=(��e�s�pM���I��5�!m�hq�8�Y���Vr�߫����k=��=@�WB�t��tG�6�$S�k&�x.c�w����ᒠ�0Lj&+��KI�q-gAI�`�t�� ��J9L<�E߬��0S��wbB���qi{�L�8��T3Ui;�`�z��03�p�x� ���XV["*4�VQi>�\.f�f�7���a���0�Eq�L���^�cLB�%*M�U}:��aX`P���wA)�E�U�dS�s u3q]8��_���'#��p,�ٛ3� �a �5�A@���"�2�Dᶂz��X5"�S��F�~��k��?LY�����p�����YO����쩱�09�}kV��#��7�J��ԉ��H�ٓ��D�v�?�Ɯ����R�!VQ���b� �iR��Þ7.����R.����{)�/�X�j�3'a�TV�s�
����}��k��e��!����~6��է�������.G @|�@ ��\N�F}����r�3栽	5b9;� z��I�˶���)#+�=Ί�ʈ9�/���(���1����(���=�e��ͦ>�m�rΦ-�]O3z�[:�뙼�jP_!����-�r*�tO��k[G�g8��8kA{����6)�N�<�-���w`4"*���)r��2N!9eH�檊����8;��l��'$cv8����Hz�+%Or-��Q����Q��:���%��$T��C�'�(�ק�c�W7T
�̋�Є%lUwOQa�Z�m|�
-���F^e�GԊ�����p���.ACm��t���~a�m6�(�k],�̯�)mPok���!8�����jN.~4�@���.;��q�7�f)���:*���Q~������Z�{Z7̏>ш=���LWS{�Ď(A[b۶�ͤ@�����P���L=K�l�r[u �y��Z�hS�EJ�D8���eǃy��V�Ժ���"���jΞ��7<8����'=���קîf�OR� ^���hb�1���8&䒐6���<�n�mЙ\�0m�Fh.��Ǖ�3��fG[�R�ccYy�9�"�{�0x���r���	�'�	`Wk�uǷ۾�3>�j�]u�9�M�hEK�աf\��gC����'��nnt�5wϹ�X5�4�����v�^�w�
S+W��cY��[�P�ve�Ǐ:���J�>��F������uv���Ғـ�+�������ݰ�;u㕪���#%�YCC�����)��������\���W��;ԕ9q�{��L{Ëg��__1�S�\5��Ym	Q��(g)�J򹦓��́�+{B]n���_��
�5���u��
ױ�!h�89���� =c ��N`���H{9;%�"�ˑ�XG�����iTz�4�A�uEjP�ӆP�_%�'ҕ�SV��h��W��Ԏ����
c��9�9�#F�v�Q}~�v��-�L`��<�2/�Ʉ����{0��UF��!�[�RS�A��8ҩ/�s��A}��0�&������
�l�c7�����(&�2���W�����*���·5)�1�'R$���h��/z���5�>�󷖐Ѵ�#�F�����rT�RJS)���Bo)-jd^�)q�1M��24�s��ӄXK�TH�{���7RK*�ʇ�4!>��o�ӞtL��V�R���kN��T��BHKL�2�G{{�3JVZ��疋LI�KF��:ܣ���ɧ�)�d�h�,���Ǩ6NP^A�ҥi;��S���-���Kj�Nߒ匨�OI�|�la�ޗ k_�k�����u���q?�5���%�����=��Ԣ���61Sfl�<���^����'�K9�2���:���9!��o%0ƕ&�N͕��o7�L���BrE6K �	��$OX������[�����~K��h�����y��u�g��]o�3�I���vY����z �,��ǋp1{��,�`4�=�!:�)��sԟ��gg��7��_;���K�+flӽ|��Ұ�u��J�%W�����M��ց��P��}�;W��J��J4j�W��U���T�g$�G�+�H&�
���E�t��y�1����1�Q�3�A����[��4puhS��)i����7u*�%7=��M��4ͭ$c����a5�[�_bT��R"��xu�(�JE)hv ��4�D�wJ`c J�/"�U��8�iU��6��t֪ǹ�F4�2��\w�P�蘟 ���R��� �6m�!��0�!�%��}Q�_�1��Ǯ_����.�uJ5���h䯢�믪����ϫ��u�R�e�/�w���zg�ޘw��T����|�o�Ŏ�o�����w���v��މ��zU�ަ*�k���_ė?�w�=�T�|��8�����۝����}�y/w�ۍ�v�ݫ�g�a�2\a��x_w���O���$4��f-z��V5�M�Ǝ�i��i��l�F�y�I��Ak�:��Q�T}�'��וL��N��a�/쇁����~(x��Y�*Y";GU��a�'�T}������;��ϻ"�w�*e�]�b,J�`QA��w���g�s<�#��P,��;�u�¢��ޫms��{엤T�]�EYn�rYF�N,ِ֕� G_؆P�`�A/q�����=���ѧv�����:`���ޤ0��[DO�Iҵ�}D��ǟ���*���a�A��������|r5{q*�bb_�c���l�1��]�N*iJ�u����o?ǋ:^��	���'F4%^�v�jΟ)�Lq�_����C'���Ҿ7�4h���H�d�?�v��⫑xP!ޠ8���(xlʑ�{���%ġPR�
��#Xy~":�Ī��ʵfL[O��ao{: 6|oL"��:�3�8�5"��N똴 ML�K8�TSO
��A����Y[TN_\U"��*-q��=x�	&l�� �\�q K��{���K{�d9r�@x?����� �3[�= SU~I�sfc���C$|��a�������)cw0.�D�d��'��_�.0�� ��C�~˝<O�O�i���E�!X_�?�Z$M���r���x"�Ew &j�K�ώy�Qv�!�Qd��ʰ9�!����'X�2��;�LF��Y��̹I����������-�($�f.fF�{����`�gټ�6�g����;�AvzU%�ط����f;��Y#�0��m��˓��WJ�+5�bJ[8d��T��͇3�r��<�2�o-��N��Wq�:����T��$ˀwѠ褜�×OV�4�$;�0���9#}�+N����<����mqY
t�~\4��	К�q�"}J�u����ΐ+�b�/roP��5��|?�}�^����u[$|f�v��%N�����5�`7�%[sG.ڗy����������`����w�y�3�X�%w�ɺ�?�s�v�>�<za��.6��89�o��|����+�~�.�����.��ؚw̉�({	��*��W�FP�VþU�U�ž�N�i_�<Gg40��K��u^�C3�/�ba��g�ڑ��ɫ.HI�x~��1���W������R R��6'�}�ns����V����u�Wgc����O/�O�F1$�S�ZcK���V;!X�Χ>�K=���gg���A�ޱ�i������{Wp��z� �{V��i�Ƞ�C/6��Bݫ�45S��B��̻~��T���U�^�l� ��C~8q޻y��\`���ҟD��>��gԌo�Ns�E�������zZm�iNևVYtg�A^u�}�S����І�?s���.>ܪK�;VQ��gZ����ٱ1E!3�9����T�E�3W�5զ�k�4�5�el^�D���)�q�d�Eo��2���Ҏ�l8$���8&t���9���0�����w�;��]��U_�2����6~}���ڵ~�49ٳ�ɓw_'(���n�fS�"��-����ϧ�(י�%^d����ߞ$������|y3�>�>g��|���0/�����D��$�5l���Lܹ�aQ��I�'�]�iz���U�挅`���(��oCMJъ�Xr}�ޏ:��|f�E�}R�U�#2�|�����?i��	��HYw�����D.*Y�h \���{$%BRhq�r�8j6D�Y;�r|�V7��v�S�$�Ձ7�@���+�*���)���`��)��Pr
M<:�S�\2�O#���`�u��kTY��Auĭ�g8<RF�!:S��bզf�pi9
O3M�O�E�������E�R��ȑ%������M�&�b�����1��Y���שY��$���`ȭy	{�EB�S�&&�-1{��OC�%�o}��� y�O!7���Ԡ(���4��x��}�C�_��4�ŧ�D�� O�ۜ�M��~�44}�y-�����s>4�>��D�55���nZ����\�YJ�=�'Y�Hf��	�W�\N�+�*W�w�T�;b9Ի=���l�H�[A��F�1�;D0�z�F��I;����$$@��.8@t�;I2�?q�9�cR6zG/U����Q�p�X�*wI.y4�O�E�ַ'��k���Wc%�pe��w���6� ��Z0��V�@��.>�.���;fϨeg<�� 9��������Z�`DEEF��ݔ=͟���6E���[褃��-XL����h'��K�˹�b��H�ˏ���"m�*G�I��hya�I�9i�V��q��E�:b�و��A�ηvJ��t2�_ww51�k���C~Ա(@�^9O��s�@a��=7�d��O�Ea��uĠ�����2�h���1��%!��us�F ���)GkǗ����&��z���X��j˓=��X{�b�l��j�)�C������|g��O*��%�HLOZ�4�A���JaE2Utb�B3�p�?�$�+/V���p����Me_t`�Nc0�U���G��K�ڴYD�i��ۻƗ�	*w�������量����*���n�kr��&���z���L��M���g>a�K�~����{M�B%�A4�p8�8r���v�!:O�-W/��X���}kΑ��}��-d�O���E�<�&������7C������o�RĂ̙3'=�F�[Gr����ן�E�sԹ����a��J�7�HCIU��/O���k�EE���Q��5��랥'����\A�ET�o�ا��WN����?Ƽu��K7�8���o1o"P,��6BS�>�D����3;JTt6xV�|�a�2�_���Ѱ[}�8��f�Y�a�0��MY����3�t�<'�6������s���{���e+�A~��?��kH��H}xߣ<�,�n^��ۡl�An<��Cy��lG�5�cS��a���C��!��+��݈���� �����!�	�Co�����֧b�q�!�����P���H�餘 m����'̟�6���GI�`��*w�'F/�
�!�!��0���<|�_� ��J��	E����AB0o	�pp������>����m��c����O9d�'�@J��\���R����1 ],�(A����vy�9��*�h�������֜.���2&o�|����=��	g����|�::����T�Eb,͈<���9߉��Y׺�4捾��Y��8݋���������A2����	�J�q���sk-m�����6
��C�ɳ^��@�����j�^��ރ'y�5��"�����A� ��8piq!?�E� �"���K]��������s���oMt�St�0�ک^�s�f��6���h���NEװi�}��Z�N��[���Y�CezRs5	�����{`E��d�fk�����!Q����>����]׃��>�eWh�ItxfQ�x�C'�6sb��>H �,����1���x ��Q\DE��w������M�d�
Ѵ����Ds(�Hw�Y�疜��"�	,^�Q_Ĩ�TG�뎤,~����hC��!7�ήR��:ƥٕ��i��H���HRx_��!7���`"�˶�K~����AH�X��Re���ǡ�������N��a��ox{($m|��C&�_4L�J��I��"�t�	��;����/����h�6����K�Ќ 鑊p���8�?H
��`���ؼ�C�ժ�� *j�Mf��)�
�?h��*=j��?k���<%�Љk���f��������Z�O�Llj���SS b���!�Le���~�2�ZC�"	Y}��� ��~��������[0u������Փm��R�0��J�〟�R�]���a"i(��=!�)���<4�х�U�U��P�x(��9�f^����g~R�~���!y���'��_�I�3����e.(9[D	 ��s?Z7����*�c̢�1o�o
h~��H��E���WX�.)U0Iߪ4ןd�qj#omm���FM9ć�J�XE��ݙ�RHř0���Q�?E�Kn��%�"+�6���B�x�D4���LuG���"-с}<�X�o'��z�VZ�)��E��)��j�J?��E�<ˇ�TO����`:��GQ�C�g$0Ł�7�3���5�ҧ�r��3�C=�?6|9��[�^���Ȟ�W����� z���^ó��Ti�r��5�}�z��8���u(T ��4U��_D
��� ��6 �}M���Vk�+����僶$��6b�В9�"γ�E��s���He�2������s�&"t�Z~�P�?��;������5!�n�YVNՕj�t�����U� �CK ���U�t�r^��Q=��mO�jf�g�5Q���5�g�4C!��gv� ԗӇT!��������!�U��DH)�=�	p�M� �R�갥�CNg���w`CX@�e�e�qo%a��(��� ��It��PG����X��N���yJ�\�k5ψ�����Iτr�.��x੔sڌ㪠�QL�Љ�G�l�Q�ۀW,$Q���B�	Ψ	��g��}Q������h�{�����Ss���d�X�>��	.B�X��e������<��Ca��cI]�n`2QM��m��F�pg(���;p��k���l��-X������@�i3y�"T�M[��c8J�F��A�,s�۟��T��,�r;�Cى��?�(~�i�tI��Ƌ��\�Y�0�o�4](t�D1̀�g	�&j�"�Rc����w����'KYc�NT+Z=@bȔ�0���K�ggY}���Q����eD:Z����/uԾ�v� �p-T���#7�)/P�>��J,eQ��/�5�E=�j��/V���~ ��Fo+�>�6��zl-.zu�h�O�'W�e����a�߈����|�l!	���H�3p�	>;��Uu�Hj�#��c�y�;A�}��`Bx�R�"R~�1u�l�:��|O��Ɠ�U� ����^<^�z�R��&1����|HA���5�ǝe,���ͨ41���ˡ���C�j���~��	�ުb[U�Vj>Ad���Ph"F�UYV��?�ٺ�k��H�>������1�
C���������ƽ������ק��M��J)��*ףʃ��6S�اnm����y�C3J-p6�5qf�%۵PhHC\���u��L�;�'2\���W��q9ð&��h�" �Hw�{
y���bFo�hxZ�S:<�\�y��g�ݜ}�aީε���H�||vQ��Q����m��4k2��{�B��
�)�����?V�\��4�U�^�3��4+��Y�i}���axdc�Y`�߻i�mq=wd����PTV�
��4�n��7�/�B�'�/ŌoZpּ��\Ɨ�C�̼}�v�>�r�,L5��2�>K�Ϛ��2�өv�ܬҴ�3�]��<Kk�b�^�З���=�lnn��X��:�̚�v���1�nmC�r�7z�rD��>8wϗͫ�6R4a��ؤA ��W8�F?�m��F;px^�ہ��1$��i$��a�%�kl$�<��z��60���>22�s�a�d�vAr#i���@��Kd� {콮���`
��!|�H~��Pc����sK7_H � ��wg��q^��,���z7l��|دIkT"�v��R�&vV�s&w3>��n&wO�j�y󗽻�U��Y_
Kt�i8��*<����э(QݐU{�%�60�n�y;>�$D����3�?�E��C<c	��aA���Z��y���%"$��ͱ�	������m�׷\]�H}>>F3a��>�1��r�8�0.勋���'L�k�<�ϡL���끍�91Ff��7c�!Բ0#Mb�*��E�1΋���u�Ϋ�;<����h�0[�
�)1�V�xD�����ԶaLղT��a':,	<�j�/��ɽ5�[��[=׆�m��i�"�U~o�E-e/y"m��Gc�h�3��?:�2[���݀��Vm������L��Y4�k^*�d�J�cu���y��j��#ơ��ȷj����ZM�RM��S��f�A 8˃w�0N<�힅��~��=o��W��[��Ű����R	G��K��/Պ_�M��Z3�^,V�ui�[���y��n�[��Ѡh��%�8��뵟��nK��[��Ϊ��l�e[C������;ϕ��s����>ӉfNs?Ȗ��P85t�`��u�rt����FڋG����|~��W�iĄͣi��b�gM�*+������G��:4�lӡy^�b�������֕1c��L\!4G��a�kcr���n��&m�4�Mz�7>;+^g��m��$3̱��V����N��]��4�	W|v� ]6�_���1�����ϢN�Av��U@�s�P�X��\�4Os��Gв��p�'\Z@e�����9�Fa��P�,
{J��O�齰y���U��7�=dş����Р�s��[��J*�d�u��g�J��n�ґt>�ծ��x�*Z�R�|��F�El_$���s?ח�s5�9#Z�gČ����GɁL3���xeio�����W9���}����qA���|��U [#y�dE#��@K-c1�zB�>Ǹ�]e��FO!��$�PCBd�`!r;�?��94��݈p��Mp%cM&�H�"Y�ޔn��ь�BE�{=����ֲ�N:�2����6�OOw�
�?ֈq�z��.έdZv�`���˨� �<���՘x�Jm?e
�/!up�r�Qo��o�8�H�SMmǵ�$WL$�(�{�f4#��v#��� �����|�U�@��!�p�5�����,ɝ�!4:.���Xo&^��TI4o㽚�5�=�
��}��_�Ϲ/;��2	��{JC7|�zRV3S��KW����%�y&յ�.�j'�+,��D!���H���Fݮ���vtB�����'���2��ecn�k��{�E7����MFZ��ú�߀|D	̏iB��S����i����M���R��O��fT�?��84���� �5/�u�#��Z��gp
>2Ɉ�N��*��iw�N;u�?	�S�7������i껞bΕg9�\w���Jdp֒3�� c�%¯5���~
ڇ����y��\�ċ��S�pj 䬏�Y0%Ҡ�b���,�ۺ��&�>G����}�8����A%�52�5GQfzO4'A�b�4t�WA���3��� �o+:�Q(��ZNT7�_·�a0 UzVH �hH�F�ˠ��)a��hSezVt���r���_�d��A+�(�)�L�����ޏv����x�=޼�T����|~7R�~]S����0�����������~>�d���nfL���@v���_WtB��%ۄ�*d�~4��D'���W�[�џ!�y��Գm�[u���l�R�C&lF��
}6#yodbG����A^��A[���7A��$��5&�Q�6A)4Fs{	��	UbBc�А���l?n:��7鹄*b_�I<e�#$�:5b��ڍ�.m�(����۹U�N)�f�}� ��k-�-� ��Z�G�����x>��t蛠��TL�ٻF�)�}Ȋ�6�ضk�����B�,K9��(���{�+�O�Zb��uE�2�i�����������c�)JҌ�2�"��q�'��Pp[)��bp���vd7[�z���L��^�	�"�<B�t�t�rj�
�rl�B%�N�}B�bܕ�V�78�z��|��:j3�[J����4��Z���]F}�}���%�R��X�����V���G`N?���7�!qG���-��ے��i��{���d�D�1�ڧl�A�"1iC�Bw�gZ �s9t��#�x���J��B�
uwL���ߠ<JB(�,GmX|�H܌Q���ޣ���l}��,�@������9��D�ݫ��ʒ_��@%��x�:A��n�IpNs�bֲb�-�fngFw�`;C2�^�]�v��i&J�Df�_�: A��\���H��;�S�r��d��`�Z���s˰0����x�V��Qk�..qy���	+1�| 0"����
-�Ә-�J��,���R{0����	q�h��%��=����B��R�/�"?�B��b�jS���a�z.Ž�i/^�����.�7���]nf�L��S�^��uƴ�u���؝� V��Zc�+�� �ŮMB2��0�4v�m|f��|6���{�$�$��I�̎AU5��t���!-s'IV�oMa��<dMg�1�P�X��,�f�q�!(i��C�����10aIl&˫�2Qlo���w�F]���ֈ}� �C�g���4Y%��!�lH:��/*
�H�j<A��%�'����m��Vpm�~�c�� [�}.t6h� �?d���_~�b9/橛�@穸;�D����n�
��	:�$m,�k��D���G̲L�F���3e���BPY�A�Z��A�����"��!�dYMj��*(������v�(Y,h@�j������<��H��!���_�Tz��="1���g�����n��c&2���3�d�x����X��,ݽ���v�~f����/1o$y}˛i�r�QPj.��H�ssM��c�l�m�}!(0x�d_�i�8
͙�����@���~��w�ܗu@m�����9L�ߘ�ː�'�S���~�oi�Ӷ�_�p��@��,��S�1�)f�<��:�!��P+A��z�P���h������s���`|H���RL�"�u�ȡ�'�/k[Ai��Vᴅ.DK�.����9��ع`>�v�Os�uT����o=VF��I?��/,�r����En�r��*�m�'u|Mj�ϙ�`��̖ws�V������en6e/OZ6��V���r5+WӋ�F �=�g���&: r��R6�O�ި��;�b2�WJvlO�@dr۔��l���M;L�)~~��o���Qw��"�H��[���/a�G7�0:p���tVQ>
��[�\���!�i@!2�̴�J�Ǡ;-h:]����Y/��l�����LѨqI�o�^��LQ�c[<T���ܧ�َ0�z�5�}6�	Q�\mL�-Ĺ.:�lo�����e�k���ܠ�����e�Ge�Oe�eY�>H�µ粮�Kй���u�42���d�幪?�,y��񭪎�����
�Ϫ֧��qY։kY�	ŜA�% �y��5�D����8!&�!� ����9��h��#� ��}1s����W�d�xk�x2�9� _\( ��/�����1@x}����;�Y|u���z�U8���x��"�����}�F��S�GZ�h������&nM��%L���B��m�:TE]�]�t�k}w�|�VgJ��@����e|Ӧ�J��k�Ny"܀� t}֔�NaJ��ڹ_�N�~������ΦP��Y6�L�U���n�8�iȐc����]�B5_\�sc�X;�S��`~��Å�u��z"%y�������-�r���/!I�$#�a��:�y�ED'��]��P���*�n�ׁ�����^�뿇7���\N��Ǵd�2�!o�{3D2�T���`�К��-m�� ����@�%M�SC��ɋk�ƥp	ء졂#@C.�I�pBQ��L�ˑ(�ݧ�cl8 ÂQ��:$�����j�҇`��%A;O��=<���*S����Ff�c��P�Pw�d���G���j�tS�1b3žG?jLS��ۦ��r`>�b��8��̩6zKyN�����qI4�Ju�*�Q��2�\��-��͓_qC��";vb(8MkJ?�N3%Wg��y���ܣ6oh3ڬЮG'��ho����ABYד�OȌo�P�g����g�,���y$���¢����R�^�5�:j��!�(�;���Uv���SI��^�/�S�2�%���5f Q��M�eu�Ά�芧�{����ඡn%�Q�}�M -�L��&��P�c�+o�Ƌe1����d�2�p�@3*�����Ҧ|/m�%5 y�qul�ڿ���6q���j����l�c�5!��R��H��;[���5�O��}]����<7��)��0�1qC-.�|���j�ӜMݶ��7�9p��`���@P�����zI�l@p7����7 oz�k_�#���2
��rǦ���Bz��p�(I �����ws��Jm�Q��׀"�� �Q�L�{H=6�j�A0���4��p �Sj�a�˜��۴���y+}	MQD��`�?t��^n���	�	����O_���s��#���w���O��6�&B��i�%���f,�yx4�Ӥ�N;��w�Q���$2E(��gB��x����a1G�KHm�����:����D>����&t��x��	�&1��7X;�ڌ����H��vt'b����@�v��NL�u�J���OQ�����Umj}Gg�j�٣*���b�Fo �i��B�#?㨽 ��,��4a>�2㨨��k���l��nQM�[ ]������� �n���{�4LD���w@��;Ə������XTs'JK�j�D�jZ<l� ���c4�M2��꼋�;ݛ��c��B��n�9?��7`d�U�vg`�Z.��L�(
����)�w��)��iD���m��ۍ�i�_&��/�ij��)�ۉ���CA����������L����Q�::\LnT�ߑ�{5��=�`���Y��^��m��y���u�\gk_"X3�FW���[��1���,`�,U}�.�.̬�,V��
�l�"�Gߍ�O��h�N�W7��Uq_��+���Y�w�����ŔI�.H�nbj���\[fڱ`���vo�92�_W~<O�z-휷8�P;օ�A�;9�{�pd���s��PW�c^�����C��H�-���JN��f�.υJ3 4��_��/��Ee1�	���=���|�h���OM߿*�+v/�P��3�f\�A������%�ezbe�5�=')^��ڀzDV�ѡT״�D�RV��O�,/���y��2�?S���Ծ�j9��W#ě֑��}�v�#�$'3��/�]T�-"��K& �S����^ԣu�SI;�߿���=j�Ԩ� �#��Kt;�?�u�L�T��T�Á�(v��b��q�xN�E!
���^���~�UK#O�=!Q�n,Tϩ�%�T�.���Y�'���\v!���P�����<���5��F ���Y�����ɴ�2=�lc� V�뼳ye�|<����(Ef�^A�����;�=l�71Eq�(U
J|��N<�P6��JUs�)���3tK�vZXS��;;^ݔ�g�������-o2�Ӡ���]�w�,Z��OB&�ǌ����t���Z�li���AH�e�ې�禄�C�+d(~ʇ��B�N�Fs~�^����6A@GDㄠ��$�N����l���L�T��_/��s<�\t�ߩOW�.�x�_��Iu�o���d�_�+�h��sAP�ZdО�C���d�d��A����n��4j0H�gFꕁ��?��Y�� X��f�?�#����ܶ��֞���C�������W�Ʌ��FZk(|]r$߮������ϕ�+_0�_��}!�\�Q1���ę�zŌ��B��æjUoM��~EQC ���͂��ԺzP�O�^�����s�!u@	T3�|�\h�2���<�E���f��brޗ�Uΐ��3j�����/����v�% �6rs:lǕK}�e��nO.�r�=�]aPl4��g_hfO���&�mAL�$S�.˨1o[��í�Ť��l)3�`��"r�x�Z����ܴ�u�\���k�[��f�i�^w!hb2��s�!��� N�~�n�l��n?BYZ{mp��H�o� �����9�_�-������SF������c�9ՠ�Z�L3�����}�L%�A;��c�A�Ie����)��Ǔ}+m=�m^��em�l�uµ��Z����ԶXm�U[��t=RL��#֘�l56vR��E���3�E.�+sz%fKP��8X��ͪ~���2���8���j����u�z�����=���xHp)]]�|r	�sΉ5L��p*;��)������[��{�tZ��@�P�f˲��P���q�26���L�bj4�c�'QK��Ѯf��=8��+T�X�Y�ʢ���T���x�@Fͫ��Y;����ݠmer;�X�\�_�����x�G5:�ZsKw���{kQJ��x�Bd�����|RK|+��`�j3�PK�d����i=�T��=�������cQ�c�2�YO��z{s�A5����@)��
��Lz&q"�n� �gt{�e��G<�osz��B�F��ϵ�/���_����,��K�p�����K�$ª�x�OI�+aQm���4�W��%��p1��/=(7@�^���V��x�v�G;��Z�ƱK��� �DP-�)�ﯴ��B�5�ʉ�=�D�g�Z�cYq�V��$������;B"˙eʉ�t�]�}I!��s0��F	����cO>fn�%�]2N�z\~��lCv�RTg-�2��[��#j�G:J�O��58��=e�M��qGn�̧kd�����Go����wXhWbu��o����WZ�a�pg��g���0�%_��y����R�����s�~�6�S��@Y��4�ϯ����L����)�n|0�a��w�/�q�T�?��|�pE�,��}瞴��#�{��co�y�'wAlb}�O����˙U�9�y���~?�~��qf]�	��v�WI"�I�'_���'/���X�]Oͮ�9�I���*�˴�j�2�����}�}��о{���P�05�W~i_����ڗo�[WV�l���2z������uo��sko�;��k�w�$�F�߽:{��Y�w���y����O��
���Aw-G�ږ��t�^d3�YJs����nB��lG���=�/�|Q����yj,,�E�ٖ2@��w����~�_>S�۰#s��:���<=�0�mʌB(Ս���h;qmE�p�yᎮσL�L{�Y~�D��4�����I-�Dz�/�m���E��J>ۆ=h,/�07Y]�6��A�����j�s�g�G"7���kO�\`"L(M5���9^^m�VD#G� �ڼ{�bLlOM4�'����^@���Ҝ(���;�N��i�ώ џmP��vf(�*��^P�A�ç�3o���B��\��	������;#Y]�,W3f3�9�y?�͛���?toG�R�����zq�Qos~kq�E������P�kHK+�\>�ф�������ۋ�[Al�MD*����_t[O2�sK�H\- D�e��<d��;Bܯ.�U�[����`�t�. �Dz�v��hp_�vG�a�.�Dv��[�p������箱�?qvG�^�	�G�e�(����4��k�1�k�`$����Qg<�?�ζ���"��"��h�D�M��o�&��2��g�G�W������E���w�q��|� �E)M��0�A	�#ɑM��G�VI����.m��z,e���>�PB��0�=S���e����DW��8�Vm�+y��z�`a�gFh�ب5��+΅�1���5r�NK�m�zS̹�M�m4 T�;�+�q�.���-�����ч_�g�V�ŻSw@-|�![e��><\��3{x1kQ�B���0O@<�(�	ޑF)���J���@i�SL��#�$#VbJ*�N�,��3���+G$L�xl�U�-�옳�2�Q��Y�.��ԭ�$���iD���>"{��T2w`�f8Z���"G�R���]�Ɯ�Kaf����o�]]�k���j�w;��L~Z=`������ٳ�M���=.T�Z�za���F�@"�Hg�g��ir�=���Z�4%�Ҵ�3���"�cwbIUV��^����е�J�<��<�gƻ�Sqwr����Ӄ�|�}�:���MJ��L:�fwM�Ω�e����*���i�gV`-�ۢ��!B�m[�(�ۜfRR	0���m��UTO1X��ӵ�f]�4���]�0)h����[ȈPA�
��C�3��I��
JvЋ&�x��B��ffM学~���k:���YFX�_h���r�����
߾��R���q,}G����"���=��=�)�W�p��5��2Zx(K
"�e;D@�Z�繈e[��֭XD��Y���\��^�8j_<��V40� �c�A7����j�3:f?�L�}�T�U����{|m4r[��������ݹ�34�ʑ�C���>ٞ,���<i Ki�ʚ�s#�
������V�M�?$ϣN�L?�Q�k�+��GN��>Í�62b�j�o�%^][HHu��ꧢ�\=O�bR���&V^�g�b�����+�E߰�,�b��$Ř��L����3���c	�~E�_g�\�䔻*�Q3�@��H�b���Ѻ��7ף[�Mu�Wp�N*��s����UJ�{��t"@_dD��c��/cg?�R��]�{�]������˷�q=bĚ�����r�d���R�s/�� � E�`�M[��Vi���)�A��x�,K�Ȣ-R���O�|��N+10o1��zg�����y�u�iiD+��[e�4����bk("Shu��۞�R:�2�|2�J"]�H$���&}(N :Vf���M��1 �e���7��� �(^�cD�NI	Y��z1�s1��6���b�b�^��E/�Q[
ĚLx��R??fi�$�uR���I����&�3�_L�,/��:��W��(�Gyv/o"a��,��Z���|
em���wle�s�M�	�U�msIh�ɠ�����+\�ҙTB�DM�vfS��*���~�nS���1�`\��\�����?<M�>C�����l��`�YW������z�vQ��+����R��;J�
�ʆ��r^������|�L2��|ϾJ|�M�̈���N�3���O��ZZ��z�SB�Pn^ݩ�/�cj�Y7f/��ݼt�PHUcCM��D���ײ'�Č�K���=�n�Rh)�����ugIeʷ�/�Q�K�p�W��3����T��cР��t��L:��q�V^�<C�R�����O�A|����tɮ�0�`(�]n�Y�P�1�-T;�E�FZ����as��ܯ���~gB:"N>���T]X+[�;�c�����p��bGW��m��̯F)�U��(���������8A3����=d`1�j��e��n�����P��M�)/�l�ͦ触h?�!��,E5|�VW�ޕ0���M�-��{j��T�z��q�zo,�1��~��bG(��
x@ (�{��a��S�G����<��h�8�J�I�8��X�y4��B��ׄ[��,�06e��S�{�Ƈ4t�s��~˰Zu&�B��*~���(#^1*,�8UV�O�Zg������~on��,���von�7wU�i��$�n��S�� ~��s��d�Z��$T8fc���I$2�����6z����&��3�.b��R*���(|�3�H(�9CZ��� ��Wt��T]i�)a����	��m�ޅ�`l��A£��kD�ڠ��@��k�r�q!�qҘa�'�* �7�l<�}���H��r(r��Q�\�g��t��O#�$�'IuV���a����������.�%T��[r��1vu2S�w��c��S�@�G2d#O�E�Ϸ9M��GF���b)g̢�v.W�x�:��7�n��IY�	�����s�:�bCxA�>+��oi��P9���s��6�3�R�=`�~^�p���ނmB�"�\(��� "�_,�]�b[�Ŀ\q���v�'<U���������.d���j�Uk'��rm��-g��!�3q�
,o��ǥ*�>z�3�5�D3�R]�Q?�y�\���Y�g3�>�4��'��+�P����!F��G��������w�;����W��-�ar.��&<�6cޒ;��$E�{��ʝE���-`r��-g:lb��݄j�uE�1e5f�J�w�aV�h��:������cBpEX��4��E��=�t\��*C*v!}�ޫl��ƞ�����Re���Q'��@�٪\uq���/@2&�pK�4�˽���cU�/g��}]��%��YA�(1	���|�)�ˋ���������;��ļ�T�I_&�Gߖ9���,]��"�HcKR�:����[�[�k6x���]��,�4����d��'*MhY@������@���nt'�9\ ��ͷ}2��T"�w��`;^֠8�)�!��U�+>J6tGG�D���ň�
H�4D�`�(�>��a��c�c;Di�4�)���	x��g��^��lì�,�h��#~E�d�� �3����E�
�Kl��NLڌV���&��n늙���ރ�w  ��+9�q�m�"8�����w����x6;υ���p��\�[�����EW������~❷��b��<�@�T� ���X�iIJWF���F�}��0��Y�NRc��n4�/�r)C�D
��f���*���b�T�;��(9�q���x�o�Tp�E��lk5��H��O~Є~יR*�����4��f����X�P:-��Q�����y�r�q�M�~4J\�q��F(@��a�n�$��؅:�T�N�B&`��8�60�jHl�0"��@�ޡ��Qa���ܡ���wl2U��!$��8U���@+����N��'f3t&4%7A/Y\W�r�?rMA��u����{����u	�c��Lu��y/�o�1��x�\����T��VҮ��I���|�����A����%}M�ё��6E�)�����ic*��5	�;��=�pug.��>���Y��e���XJs��Q�Ev�:�TB ��p�Ie��PVD@�1��,u��柨9�(��Bm�7���a�˴� �\��AZ��1T�Y������#6��~�C�����̓����
�(5�nc����`Ao?����j)�D�~����6~��̠։LhL���]�q9u�SZ?6���������,�_�'pHkP��^IM%�~��KfF�2O��L21�!����C���^�:c��ǧt�K���i�Pԏ�g�|�5�#����e���x>t�rL�����v��J��$��%u��}Vb�:ƴYy'9+)�Ym�:1󀓛��8���:A�K>�߷�d)�����Qu�i/�}X�gL�'����E��B�v$<G�,;�i���^©]�O�~��� ЌK�ч��k����?��<���\)���[%~�������$��0*�p!��_�)�sL�=\� �a� �(X�HW?�=�}�v���ӛhp��P�Z�<�6�@ꥣ~BO!1�Dd�Ρ:�?�J�0MX:�x�(����(��{h�׍?�`G�8��m�Fzg.�Tt!�+(:��#����Y��!ǝ�*s�ޟ��l�&z�3o�=y��v>�H*�Y����MEY����,3UAhx�T��q�*�}e���/�_�����O��"�+��F��ˌ��t�{��*�4��uqc�o��_{|{e�ۧsQ�i��Wvq�q!��Y��9$�6�<n��� ��$�RO�| ���*7�ga�鳘��'~���Uli�G�񨇤Q�G�?^Ǉ7f�����8?��Sף���4�����S�E40U�v�*V3&v[�+��t�i5?t�<���aE����<#�蟭5T��[j�iA�C>hs�b6��.�1��jR��y�*�	&�����PCA��� �vwS,�<�*�X0Q���"9�,�6 )�:���;:�Wl
�I�ﺥE1�6,h�y�W��ZV��I3�5pb����X�c�W��߂*���EIv���"��`�2�`��q�����\X��qV��%���;�3`�O>��+vbG屭��M����~˪"ϐG�����R�{&��w��ьu]c�ƺ�J%՗ϒ�Yp��9������/��|�e�\�S.��^]�ǟ#����6ҳk6x+��K��?�Y��m���q�2�gB�3�Sj�_����<N��F�nY�� ��9x}���vY���gY��f~(�wU���\AI5����a�y�E[����T����nVI�uQ�/[�|8�hTގ 2g�S�j�bmK�:|⸤nQd�R`ڛ��uq��q&��x?(�R�6q�na�0��X��-��P�\�1���+3������s��A]�.TU�9{=��1����P_Z�`���.fZ������V&�X�wU}=�p�^��>\���-m3�����x>��Z>�T�X=4˧._�鏼�G�;��;��jP}9�ˀ�J/	�AZ��$�j��ݡ�h��AL��)���򰃢���=ʂ�����?֫�:���;
%�~�3矃� ��Z�D�q�Q� ���r���0���=�ksHh�4 ��ө#��	~Ec%�Ry����u��c�c=gЇ�9�&R׿B9="}>�$d׽�P�Q��v���m'�����8��ڧcnqݵ�+�!�n��0�nr�Z���g-���W���Փ��+/߄a�Pfy�2k���y:����kw��^D���R�"}�zP/�+3����
�odͫ�_ܩ�6N��Y<6�5yevӁ�����kz~���o^c�}r�l�p[Sl�P�}K���֙�B�$o���o\ﵵ��pϭ;\��R�7��>�W��͋������������b�&�s���Gw����X�{�MO��{KN�kׯ��d^$��dxީ!� �'Ɓenh�-(�Q"���z�<�c��/A �ִm��=b+��놃;P"��� (���!h�,@���Iֻ��¢�M�Z���C�����`�����	 W�=T��$m�;�V�O�����fjrmw�:�{�m��l�n�X�kg5�zT��`��6�,�Šu��K`���s�~:V� @�б�$��w1��!GڅĨ��yΌ�*t�C11�{;��RO-՛��)S�AAŴ<�#�hFP.�G�
�܆�V2�drg�g���/�'@S��8�E�?NZ<���^QP\c���&JZG_�(i]R��əgڴ�j�4ш|@ԎA��u4��g����*Z�B($=P���"���R��hnX����L;
�O@�ͼW���X�/��O���w
���|	��a':�R�%Y��i�8�y�蒢��0m��p�"��RE���J��ʁ�=#���ن�݆�	�6�
�Jz? �ZQ���e��3�VlU�%[a��w�vr6w�(0F7&��i᱁�1��O6�Y�5䴾=��ށ�$�6g��X�� V�l��2n�	k7=i��~����.�R�X��>�y���X�ys6�.K�3]J����h�dU�lȫ�ɭ{�پ\���R�6��`���]��;�T�@���|{.g*�>7�H�{��)�R��k��_�T�9�ӝ �7ꏪ�U��UV�,K[eQ/ˎ�i�����1g��T*m�Tx�����\���+V�~� �3��ޢ�Ѣ�Ң~�"�L�&
��%)$�-�b��m*�n\�U��Ӣ�?�J��C�4I�=�Z�A�P�xu;z���]��.yܴo��(�>����>�?��G=Z*�; %�o��= ȁ��
�Ӎ��+��E[�G�13��\���^4[���m��N[�BV�	S�[4�wV�f�ϘdT@4j�RŤ�V��%���K+�	�pV,���T��8�K^v�Yl�����4�J���㙤�"V������3��RaE�'O��F�٦ ��(p+lѡ��6����Ĕ��s�c�z�w���b1eI{�t"ƷY�r��pt�؆!�L�g(&|(�6CY�����E%�o�GT	��R�{ϛ�<�L]T�g�:��;���6�0��>��BO"f ��.⍎�v��Ȃ����d��������-.���4|}_e
)����Z��$ B������Vo���m\��D�B��u��b��e:%�p�?G�v���`��9S&i?6��o�)��O�SkS/�ez�"t��D$Ӯz�L�1ɞ��b$0�wCU�ZD�T��"Q�S�=�Մ�g�s���K��>�}�:�)�n��J���JU��3醋��D��k�F�;�D|9jE�r(�J���X�GO�,�'6�t�Hl��?��&&!f�~}?��9S�ˊL#+UҰ��ɦr��VL}�{����3�V��$�I;�^��K!�J
N�e������Bm���R6��rƔp�!���]�	U>�	�V�FWD������z�[һ�4��T����1|k~,:�#����Vt��>���9(�ͥ\UuP\����K�!0a�˪��DQ�PrF_�Ҍ�G��{+(xE�P�>��P���r3�c&�4�`��YhRG^�*ߐE�]���/c�ɀ1&���r����mM�Gh)G���R�~}g���9�MEГ"�D��tT{hg�Q.� �GH$��(C}$gmRn�(�ҫ!-Y��1s�����/��X��yj<��D?qx�����B�ib�%�O�_4�.���Vʟ4W�l��6�,P��S�<ĕ�Ue�1I�­�2&I�;�}ДS����G�HB��C8�K�ڟ������1�=������L^�F���\'c&矔��sل��,Օr7�S�nl	�Щ�u�p�4=fY�M��֟��Z׃���8��*v�XB�5�(8o���ݾ�b�J[H�X'�*B�J��������>�ܱ4\��&@4�</�T0�ù$�o3��Ҏ��Ƞ���:�4S)�����f�� ��t�Vf���i`T��?��K	��p��V~��tU2���Z8���~IwK_80���T\�"M��W� ��(�B*��ԃ�"�Z���R,�7���
нČ�K*�S�v�x.R����g*�-���8m@ ��̥��Yh�a����p�~��1$������0f#���
,�z�:�.�jے�y�>��IwSB!��D��I���a4�\�������/�v��1���X$(Dx���d��e ����͝�D�<5�4����ǝ���\.Q�;� ��L\"�!R�xJG{���	�f�av����!�������x�s˅^$�]�@76¢Rf�a�3i�d�P������`J9Ֆ��\���[��O��bNUy�i�'T�J�1��t]�o�����Z����R�\���Uتg���S*=V2T����ɊY���k>�g�Q���8�7�>%Wo�7��8���񎭺�`��8L	�gP��F訫z�qέ��ӻ� 3��௖
�E�@S�� *_�2�!��WIr#I��+��b�����0�@$%��T�͡�*K2V_&���a'�^�"��9h�W��+��D2�N[�}`�pEJ�E��L�_��k���:�� �&�y�i����T��j�v$B!����\���f<��g'�4)��F(� ��8鈥Ӈi`C�\�>b�UC�vmL���AHp:FĻ�_m,�q�f�#^@AM��MF�vC��p�'��Oo��P$9DI����Rd�^�G��0�
��=1��l.���E�����ad۠'�#X���z�T1.�T�^րȊȏL��'zr��m�â[<��=hև4�J*1���Nyk������%>����$ u��P�(��A��$�GR�--l0��o���Q�׶��L�Ĵy=Yg6H3B�V��rgކ��EW)k��oY��Ì��\6�ˤ=C/7�t'dKDݐ���Ywu����'�e"u'�i�8f�W�J*`t�d��,:w���M�H��i�]��[�ϙa���H���usi���2zaF����Ĕ_�Ż$���;��G��-Kg�h�b�����v�����A�$g��5�� �B�,
�	�Fʋ%5��
�'X�Z5`�1kJ�då;̅�A�3^F�#r�F���b�8PE�u�%��t�������JJS3'^�E6�"�&��|ߩ�(��o=�6,����AS��A+�ՃQ7t���3�Ɖ��)}����9�<Ѐ��~�ζ2z����X���q�YN�<�1&]������4��my ���-P�@�n��mm�~�4Q�r�)���r}���0
d�א�B�@@]�\_������	��0�:8�4��,��	�"�!l�Z��y,���b�d������ލ�c�\�4yZG�S�N�EO�S���/��t��\ώ5��t�X<�1�4��� Gt?1#H�H����)$x:Q@����	��b�$Gݪ����F�n�W�,�K��
�Q��1e҈!! =���MK�����VV��ܦ�u�n��Q<�2�-Yz�T�P؀74��0\�z��{i6i1�rn}��*�|wC�A�CZ,\&�h�����j��#
���3Y�G0���d1�o~e�j��h�B��:�^b@	6��h,[������C����k��M��ME��W�S�c0j���5�|�f�� ���	���	텊l�-�)��
���� t�i��*�'+GoM���&��;b�
��Kx�����'y�카��<���8��ʃ�):�*��q������'�v��O��W+F��t/~�i��ʱH%)��R�_:��{��тn��"%�霜-�$%M�h+$��[�ţ�S��-"�#�yܤ寕m��$\]C�υ�s-�TE��H-�n̜=]�|F���q>�8����1*�s V����w^z����ފ^i���0Q��7�^�-i�w��M}������uU�yA�f�V��ȴn��ʇ��:���@y��Jt�3��=bB��'��Q�������
�OF��eQ���ߛx�H��Z�=��5���8R�
�}�j���?|��|w�ԡk�z�\N��H}_F�����ɨ�܌�_K�pc�+��U�����G_q������}]�}V���ps#k  NcG�z��da����}� HAI�ǽ��7U)�� `�7�{�>��U��	e�F*H%N�:H�#H��(��!��+6�K�>e���g�?�~6*�����a�;x��f0�?�����mX��i������a�4ﲷK9f�ܹH�E����Ѫ7S1��R��]!r5��?�s�Gͳb�yF�j~�YQaL��%���aAV ����{����E 峦�p���Rbzs��;x)���f���L7�t�����Uc�zވ�j6*���9��lz�^��S���|�;U�x����b�HI=��_΂�O������n��rɈM�7�g<� �t'��_�<�� �..�ޒ�S��k���n��/G���i�Z�*ˆ��|KE���T��c��ţM�Y��T*��D�.ͭ���>:qN�g���oY�����������AO�� JʫH���Ƽk�Z���kL�~���֬�<�~[)!����>�-��dx����dIS�s��^k�$$V�9�pԃ@�fx"�u�s%/Q���� jG{Ľ���zyv4Xe�6����uy�ܮ0�V.Ŀ��_d��g��OLӻ0A�k�� B���e��j:C�;*���RSy��/��&4d�֙�	dJ.�pv�
�w,�G�s}Dd�C$����;�cN�H�	�d��չ~��U�F�U�g\!Y���L��2�3V�`1���ԧ4ӢJm���3f�J]�P-؁PvwLr�	=�n!��#��5��;}�d�j�7�In�OQ�_П�����?��LQ�f�9_ׁh�r�@��'� RQ�k������I��=�x9D��å��A�����.��!}_�������3��9D�����n�Cq��y�VBdd]�֫��&�U&�!�b�-���S�������c���x��ԓ/�N�a��!)��/ �����r�s&�
.�\>��{�u�뚍/9���B���u�lR��eC�1�n}m ��wCк|o�;f����د�^���<gG�+�Jw�{�P^�2	��A���M�q�^!h%�`�"8B#�)EL��2�ͬj�9�c7��Mh�E��	�F�W4f�j����#*l�L���u�ș�&�`������}?�����՝��O��2�H{�j�ڻ�xM���5��A\O0�f��%�K�~A��tTO��u�����*����c��(��n��x-&An(f��<_��L����J���+����>���ӂNp�����'���%��ݟ��c�p��ٜ��������������n#+T@l��,�T8;�gZU���������e��5���Ͼ���O�F(�C.�O �%�'3�x0��6�� ���^eY��8�*���q��g��� �j���D���]�r�Xc!�֐P�A��I}���oǨV���fl_˸,�у���8��}�Z�S�/��yt!M�(��i�蛖�p�X�u�	B�eS��]!�p�Lg8�1W�p�|3C-���`8h�@,\���u���P�X� X��F���ko����m�w��J64���^L���{u,�g��¸�q����[Y=ˊ��K#E�Q�絑9�W�����v�
�c[@h(��X��y��"ߩ��W�1;	+����lYO4�!��㑶��,��]4��=��%50�����j:��&�(���k`b<��Œ{���4Ku��nr%���i��s/�p��4�T�Kr�=JM;BR!/���/�q&�D�-f�n��ml^*4�筄�@DB�wL�O�fN���U�Ki��ٸֿ��i�0�����n@ }ԣyL�W�*�l�L{�j�	��%��-�i*--bcjY�Ƅ������G�Ӑ��}�r�����Ӣ�O�j j���j��� R�� �C�n�¦9�z�B������C���TN	|�Es�j�X���*چ�>J�v��>��W�l�����fہ���&�d\��Ԇ�Lt4ൔ����7"���y~����ك��e-���0ِ�^�MR0u^�����З�D�#h��������Hr�d�<z�h�"��ܥ��n�RZ1���iRiĥJb�"6z�D�`��F\��z�ߑ��J�����0%�"����(P����f5�*���Q��� �3���`Oq��9���ž���V:إ�{�N�u�zc�a��F�A�NJΈ(��2-lg�bQy�&q�OsЩ"v�4�����B��yS�%Z�(sh�&>`&CRmOr\`B���B{.��c�Z"8s9B��	-X��� �X�{D���o�*W_��x+Ô�wM9t�y�	o����{�`��Aˬ4\iJ���yp{DzG�A�l�R�JB�$�iՏj}d�mjL��㚹g�xI�����V�}qLPvpLόp�W���� X��tMW�ɇ(4i����1a����(tk�m��c��+b����R�2�G>�x�f���țK�ǯ%x������.�Z��6Q������T�]�I��*�$�����h'�_����G�QC��~̼H*�����L��&U?$�hjۺ�*�xh���p�����Ɖ�\�X���^���CĨ>��^??k֦���y��7�"� C�H�囝��>iM`T����|r:�����b��OHt�e��-�x�Z�q��P�)��RԐ:�Ξ�%��ט��4����C�o3	�i��V+n�{l:�HQ�#�R���4����?OR�I���>����@4&��_l&
�r!�+�q�J�z��fQMy�&�|(��I�'zi�m}J�������_��ʮ�c
.Ń1BɱE�լ'�\�&��a�mB�t}K�݃H��̤z'�EBE6�sP�a�:z���Б������[�d���laE0��� q�jOD�v����gDͲ0��Qw�^�Z�~��(���֦�i�o	Q�"�䂀�h�u�8������J<�����7\:������K,^S��)�G��)]B�!]�z$��ی'�L����e�w�&��lF���x�FM��y����$Y:������z��y.�� ^��MU�OBt���x�U��h�B�I�������W������	:=�#ԉ����f"�gw({p��,>��W��m�ԓ(���1��|�*�4�����71l�炀_H/O�aV��eU�-�:eOkKC�������>�l띆���y�P[&s@�V��]�is�	~�~�����:�F_��cN�64��u��s�0Ahb]y����o��f�WT%"2}o�W�P�b�j�w*���G.���eM�OH:4&� z����)v"xPz�Vr&c�{,Qv�
,�e������q�2��$l0�	-{`�)/�`�����}N0�=V�%�7�)�}�̚�~PE�r���=�4��FU��##yr�շa�T;�o�������Q��{�%qt��X�&?�P"1�>�����|=`��mF�$�^L=ھt��=tL���i��v�ȋ��Γ̊H�����\�	$���,)����hp/���j��A���BM�B���>�6�3j����g ��N,&��-���]��ҷС(I���:*��m(K>AD���!�꧗�gP���V�^qrmr��u� ��̼�r����Ĥm/r[V@�giVGұ�k3˺허�������X�=���i 3�fL��$��xJ!@�a��3���Q�m�'����J��(�W8����M[��?���ٷ��s~�G��bO�Eۑ�e$̬'m�\�G���.��
p08M삋Yt[��n�[s0`Q5p��^�>`Z�7�2�L���+PbF,-����f(Fhw���$`�h�M]���\�RM�x�k*��͵3��#� ��tB:��H�
�� +�I�m��V2!�1�r q��Y�o��E��t��"Q�\ _V�R�I���FD�s�t[����2�c��Wx�bIUm�bF ���J�X�S6���q��T1>ʌ��3
�w��[���l�A.h�޽�|f�-f)ޅ��B�� aT���5�)���d)T��%��8 ���Q�i��~� "�Ċ*��4�J2���J=����5�������Q��Y��FCU��5��P#
����<g=���q�#��M��Q�hD(�k��$�L�������MW.`��A���%d���+�U3.6��^Sr��M�J��%"~�d�G�a5��d�"�@�ƞߒI�PX�1J�P<(nY���|3n�_�&��=1�� ��@�5�[ 
bn�Q��о}\E�u�ځ�DΌ�����>�������Ye�/�g��dA�)rL���W[�b+�JM@0�;�9ܽ��-GcU����!���6��Y?� �T��Z0�4���eevƫ_sq��qX��R6+1&f���J>��~�ߒ=�z5R~?n���f��%*��h�eR�)���[�c��>'0�J1.��K����p�ҲoR��c?T_����/yf�H%mcޘH����w��q����i}mX�F-ԋ�h�1D2��@�J�Jp��P�ԏ}��Y��|& ^9cњ]��R$$:S����m�bg��:3"�+Q.��X�b���y��t�\'B��	_gE�X%��Do�6�{8^�v�cH���Y���	��G%l��p	��	vw���Anu4
���YĿ�ģ+T*Oڭ�WjT[��t�F�"����ы��d�ir�ئ!�?/K��At+��0&��]���21�d�-$N��?�)��Ķ4�}|�֘��xF�s�juZ/ǹCu~�v�"~�I^v�B�`��w�et-�p�^��#��O��X���4y�d��fIn���V�*Q�z(�7:�o�?j��:����0��X���^�?FM\� �}�f;w�!�]�P�EM5n�����bi0猙�Dx b��.$�Sh��2䠮���r5���'=�	l���7�BR�6��{ضp�L50�V�=���vi1���kHܾ������*k?�׬�A�a����P!��j�0P~I�k�Ku��ֹ�����|�y_�oED|�h����l�:��Vc�.��P�^�����z�z&mTQ��\�ܞ�<�����-�yg�\{ �R�L�M��5�bh��.�6T�R]&�f�"�D����͊r�&pPc챍Grx ڐ���!{��]�p��-�j���>�ߊm�@�0,��Qs���N�ۋ��F��y�T��׭�R��%S��P�3��:��쯘��s$f��9��koˣ��ˡ�$�u����_�V���uA �T�M[�طb���F�2�Ϙ��ߩlm�9�#ا[�=�ôP���| h=uB��@P�����7� �g�a�=ѝ�Br=A3f���%�[I_��O��6`����:t��9ˍ�*��m��>SNmM�@ݦ��AM���rH�k��Y �Q��z�YԨ��S�t�^��{tY�O6�����*����:+�*_O��9��m��zO����'d��c�ř�|J��|�> ��5��2ɯ���Ц�����Q��#t��i.�T�峠��L��#1�j�Ww|��Y'*}u��x]�y�lNWu)��;ݓ�������r
pW��8'?%$�	�&��7EQ�"V=K�XN��£�}�V>�e>����`�� `c<CCo�|��֖W+v�鉖���ő��Geo�a�����{E�W<'�n,4#$��G��G��goD�G�k!�����(�o�cߐ'���3�8Yc�lhƶ۫�_��b���`?T�����Ѷ�?���
g�b�G������/j;Lˤ��T�'�oC-��#!n�P�l���2�wL�8譼/4º�Z'��P%?uNRo����C��l+nK��#q��Թ�S�Wlwq������~9-i=G�'6)��e�CeGB	`& ��	N%? {�?.Y1!���}-�$We/C�2l��w�)K�����cIwÂ���XQ�Bh7BQ���V�� ��8uU�3`�L
��Z*��f��v�p�	�yM�Mn>��Z**W�ퟠ +�?v�D]��×37���q&n08x/]�T�_�ޢ�b���)�=�A�%�M���]LԘ_��MȎ�w+�������cn&���s�7�R]�������̝v��9Kl��p��G5����C�\��jT�x{�<��>US��`#������{�������,)l��tHw�S�}��x��]��q���d�5��.���(Ka�%�jw)�qy�a�ٌDaQ��� ����Te1��� L;��^�u�8�����؉0h�4�邱��0�0��I�4������lQ��Y�-�Xݩy�<O+bͫ�͟��d�-�ZǵIti�/�W�n��6X�<
�/
;VaM�m�	|����2I��� b��?H�m� m�|�߁�ྀ�¿Ou��� 
d*!wWM��n�W�mзh�X���@���
�;潅��6\� h1���p�����2��Q�w1w�fTY=�Zې��ԚFp������R[�⇯�<J�` *��=�/{k�Q��z:�&�K�*�s��yCS�\�c�B�0���b�dg�N�d�2eP@��1�t?������f%q߀���m�.��y�b��F#ï�Bk�}��Q9{K�>��^�6{���Y�\�k�e2��)�ٔ�N��*��՘Z�ˎ��8�"�a�]l^Ć���9��̴م4P�Dc�$�D�D��������ü^ܽ^tq�ʶKY�L�侱�H�g���9�<R���RbFƘ�>��H��g2�j��i?1=
�����-��:ЙK��6*8yqY�
>�3�A�:A�����g9��tS$[Z
f�O��fڽbS�k�C-�ۼ3�=��E������3/�tb(�5(T8�He�5 �I�8�CX�6�%�w��U��)�T�u_Y�@�Z��/��q��
<TV��$�k/Hvb�v��1,>`$�EX��3v �6_��%v�ڲ=��DE3��a�F�J/WI�lX���l��e�|xB�C]g� m� ]IX.�L@/���7QR�y��\|Z�k4�����a#�RM��G���w�u��;@�	,�Bԕ�WmQ��e��;h�:)�Q�L��u�}�W����p��s���t����O�'�9G�C�Tliq'�{�tZ�Jm�&�e�0:���ҫ�FnKO��յ��T�_�XZ����jJ��jy������-�Њ�����cr��\�]r�� ��'w^�_&ב\���y[�+����/�=�A�H��Ɵ%7	���j�p��^i��8��)|��3۹�z�$p:�
��jzQ�]U���_��f�DpJ�����r��x���$� ���r���CX1e��3lZjc`�&HFy=��>M���c�L)���hi�Q����waW�-���V�`oDM�%��)(3����J�W$0y|��ݖ����]����������������3�=Ĉ�u]~����.L&�w\c�?�s����u�]�����^��870m۝{Q���2U�$�qUS}�'�DYbd�rޥ;yVd�q>R�9����HO/��b�-u��hO�����Y޻�6/����g����p��C��]�&ox8VC�����o�稥c��K�3j��Vp��]��7���&Du�F�Lw\.,����~ڡH�lq����=Y���Ч;�4���nps��"���o�D����5�������6/���n�!���6�M�}��}����f��o�!WWn�:\�C�?%ŭif1������#
�%�G��;}k��E9bz�,f���I�R��ι��#b�Ӯ�m��U������)�+��WU����w�JV��V��6��(�HD�٪�d�+xK����N��e��e8�Ph�Y��M�ɱȶ�0�L�o�3w���x:�[?�a�GVH��ց�C��>�4�5$��	I+��"\����E�O���J@�uc	�M�ȫ�S�"B1�D�xd�ǎ�Ʃ4�i}*% ϩK�S3C.Y�0�����>LZ yR@>� 8̯T�p��t���&��M�&����KV�SlQSꇬl[����DZ�3x7�����w{�p/j��Z���Q�o�T�.��S�/�U�(;hKp�.��m0G���5��2���;�׻�?"p<�/
�ۇ*���{[b�����<�N��m���W�!�%%��8�Zb��!��N�|#h׺��"�6`,�C?���(�CGrQ��D� �'Py]$��hF�J��lE���RT;Ƅ���$$�ox�B���ʶ�g^g"N�X��7��3q�y�u˽S���.Afk\�u�f{���g��}��(��x�:CLj[8'�2�Mc�h�	)8V'g��R�3��?��PסY�C(���Y��S�[Fq�@FǦƹ>
���ķӌ�����d����$M�x��P�:#��n��_!y�V\'gj��χ��^B0�J�q��~� �XU�+*���}Q^\QZ@���f��slǋx-��j��|�d�Ȋi�,�yø���L��k����?�V۩��RE���x�_�+Y���#Z�+�{*��E	����m��.j�)���+�����T���3�w�RTsi4<xч"���5����Wp�/�C����9��Of��S5[�&c�sޏ�qB�a"�T������;�?&+��dD�iD�A��l��ӵ�Y��h����i��n�Ľ��#����C��I@*�F}[�&���Q ��[�O��X�J�O��_�]�$�^(�y�q~���Q��b���pS�^���9�ef�6ɫx�k_L��X�Ο��]�����;�azs��\��r���קҜ9��TaD�k)��������W��F��nr	W�����}e��jf˺9VN�Un
􍝣��d�#�b����u䏍A�=d#���R�z�+U���ô�r#�a�l5�����Xo��K��?�����bI���6c�������x�P���������3��9j���z+�dc��D�����g�#����h�)*  �F=��]�;?z���brX��� ��d8	��-iK�6�~�k��S'H�9=��{�F���A-$ef�-`�vU�&ZV	�a� lk��<Fz�J���tI�?^�6-ޚ`U�m�ê"���M�Ē�E-m���g�b6��
n/��b#� v��aeJSji v�lϲ��h9//[�P/rY.[��-#ކ�τM'�&#���ʑ��H��D��D�c��/,Ofo����L�]7d_�Gme�I��g3����,��
���t=�~�����e�O"4xgo����m!"�d��Fh<x��� �T"��K���K��钰�~���y)���v��e��k�>볪�����	[^Q�XJ�5|��+�.�(�-`EJyi���j��m����I�sS������f5I����� lr[q���\{4�{3x�0�I��l���E��z�P�YZbKFR��x*W	YB��vYI��d����K?�'ʮ'�L�*�Ǌ���P6�(���� "�z��������Y�J�ݪg�
�̋i�b6�#��J��u~�0�(f&ѯW��Z٦b��9�8�%�[�~��		fր-��� mC����������({S�r���bOG?^��䜶t99�S����
�lZ��t�%h�/�L��%�ڌ��$��l�Hxr\�v�Am_{$~�u4~^��g�F�c�I+́�s-N��,����X;M��k�>a�a��d�|� 0>.���X���~��֗`Ȓ��h��kV����ef��'	z�u�O�=��y�B��>��
cC"ʺFy�Oî` %3�x��q[���=��u�B0��	�N���.��et��rM�,�d�h�ľ���Ԉ�)�Q�Y�j��隷��(z�Z��A2y�<��%b��I�%�V��:�;�w�
�i 7+p��?����yT3nA�hY)WQQ�����p��[蓓�����'�6n���p�����O��Gi���r�sp��jǼ�KO�I����$n�&���F�J���a��WF#:3n-Ɠ4 |e�ء�'L�N?��g~�с��0�8���K�#ؚR����{����O���:���T��}r�E(�,וL���M����vy��j����i�6}���VW�ƺ|���UT'���.�'č��+�T��ۗ|`@��^����Iop۵��5�#c�/$4�+��/Q�]D8/�S/K@���:��e�ZoP�*��F��m����=�J:w7��r�F��Dܞ��e�)S9P\�p��7���QL|؅�:�s�|$��H`�У�c�Zv$�m��_Q?PcQJ:�����0�Y_�`��MFP��ݕ�ճ�z��J��#"X�^��(��o��p����M}Z�/��ඔW�M�Z�~��	I�TZ@�O�Ly�WD���%_7�������g��x��fcӶ�/��~�D�aN��_�x�N��E�w	xy�c����Q���+U���Apkn�m9���������j�-���;��7�G�A��yr�s�ȼq}M�FS[z�#K�rgS���p̲�{R��m�{�z�aϋ�}Ƹ{>:9�e�wP����ԣx_a�3���;#y�<Lwt�f����c�o{�F���Y%�!R��Ȱ+�4��H����m�M<�C��ʯ�j+��c.nk�娦`>Y��ݑ�7���y�@�ûS�E�����:m".�p1�;�8�����յ��spm�0[�S�L�Tknm�==���l��@)+!�?:�-Hc�:��n5���f���\���X�<�K��&I��i�品��SkH��,�#F�j��Ӆ�)�t������jVl��=#gǨ�<��<��_��K���a�n����h&�?ޜx�)�����̓JH�� ���`]��U�L��TN��	c:ze�F�۔6������Z+��&��*�ۂ��Vҹ[���*�*���f5|�U����Jg��-F���LB�oQ��J]��n������4j[�/��I����s��g)m��p�ߐ�>��;I� �=U���'i���֥7N�~C�PL��ȿ����O+��}�]+�f�ԱH�jd�B�م�9�Y��Z-�ٝ��{v(��Zyd�W�M��~���O�}�w��Ju�5�z�,�ĩ,#��0���Y+��tĒ�2�xĉ-��e���C�Y	��j�٭�켆Ƨ���"���e��׵�(�k['�s��@D[����#�-��^���f�*zQڻ��d�vvs	X9�A��"vS�*�i���E3 �Zftp&�� H����F+����\b�׋���e�o���Lȕ�	�I���`a�҄f���jy
����c�5�H��I.2y�����#\J*�K��I�Rj 	��F���B����b���1�F�&)z$"(t,�J�d��-�\�/� �۱U7��T=P��6]\���j�:��Yag�
�䨽Y�S������맹,_�W�PD/�z�%� �G�>�ON��Y�V�����I!m|X�^ S��]Խ���AQ�R#�9!���d2*�W���X�H��U����+�kU��fz��?��yl��L�NZo�5��؟�<@�4��SP�y�f�ʀ���=�G�������T�0�-�v�%��/AY�gXV��l5�5��L�5���)�����=����$z}��XV�b�<`���,���Xf�]CZ[�ڴ�i��a����TM�Ð�7gH�;�s���\)�b@�L>\�V����Ȩ�bc��K+��2�Y��`��c̯�nѯ0�0��A���nA<Jf� ���~��#��i���u6`)�K�8�$�A+[|OqXd3jZ�ܖX��(��(�_��%$''�1z���(Jo�{��$s���J�<�oq��ۅU�V
�v��9=���s��ߎ�PB=�fH�u4s'�ј�?`���i�BD3�ŘPi������2�R�=f;g�/k���D:w]���O�J�1A'U�a]�fI/�(E�d�%bX߈T�hXPl!H�u?�Q���"$�#d~��5C-I/7NS�G�g�R��aJ��ee}&lD(������f��Ղ.��@mo�x����E	�f���q�����dR�o;�qzK��pf�.��a�٧��F�tr)�:B�=�&ʉ7Hugii;k���Fc��=�;�-2(�����{�BtU�&[���{����゘v[>L!L�oYD�Rb����P��-�ZCzT�Z��;�wm���F(z̾ofYf�8���^қK0�=F,9�j'�"�uu0A}q%.L�F,z�xn�V�]k�)9��۽�Z�A�Qwi1��KA	e��<�^��RB����.)X��E�f�|I��u�]T��]$�����xE�ϛ��������� ���N-~��Rc?��Hd�K�+�Ac�v��v��|Ac�x��TW��i�f\��ku'�𬺢[�b-_�5�Xӯ��/k�y�jm�Ֆ`�� ��Zz�I5�Z�o{4r�T���V�G���C���v"�ڙT��N6�\�U;�ڜ���b�o� ���@�Hv��QKc��ւ��I,!\��KJ����|�:&)��q�4����7�"/��;� T��)�^��Qo!it�4�ѳ���I�Ű����c��$o��A�����:D�*sU���Z�o��.p��� ޚ 13U�＀��3z�n��ވA�U�8Ӌ��QB�;�o��ǳ;>b%��1���!����8�ᘫO�a�Z�'h'-��Y���>Sl�-��P���F����_�Q���v�Z2SĞ��$̇��v�>��>��m��P���E���:���xT `���ΖGcy�e�EѠT[�m��X�w��'</]IYn|�8���D��`T�����m�T7�XXI:)=�#�)�C�!�3V@�������ZLZ�1�-�F�;#�M>f�OC��!�l�i���#�mz݇~��з���}{!��4��2�u�������/��t�����f4�I\�Z�7�����ߛ���o��g���vh��韚4��eg�Z���ӵ�I��Kq,�)ZC"�����o����1@#r�˻+��+��V�����T�� ���5��
C��K�C��	�OmV�g�5�B�Ț�%&�E�8� zx[���yع�!:6S|D�;ׄ�ʦ��0
ʎ����;�[^5Jh��sy`/�>C��3ߜ'5�cjLz��z;bV ��CJ���*I�ׁ�>�/�$8��6Q�_7�L@��g�G��
~b�A��`�����c����8B�GH�׸����6����M�	� �qoD��`gY��OK?�lC�l���_��W�v\��&�ȉ��ҌC �s?��jN+d�,q�yBG���Rul�F����]�v�U8/��BYc���2~�����&8R�}�K�+Pl:�j+�EM�_��D�8��&�ђ���t�۞A( �~��|g��9�/JP_!�JO�j�^W��u��WR�
K\CU����9̄�lh�J�B3�%�̇����������� ��SH��ECk\$�j8�.�����w2��B;��@��'�����Q;�����;W��%�\J��W� 9��� �CK ��!�