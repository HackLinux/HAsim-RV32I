2�]�Z:h}�8�
���j�����Z9�^�%L��FzZtZ]���� �6z�"�et\nib_�����H:���y����!%�dB�[8��W_v3�8��M|�?ά`�WU�3}�~�aA�8�#�8�Mȫ�:x�S����Gmx�Ko��7���fő�-��r���Y �;��e�L+��, F��6+/��.�{bL0��hiY��by��?�B����7��=�֏3|�͢2������>H����i 
2���.� �3sW�&�8�v'zm�}:#�2R�'x7�އH���Q�K؈����?�����ά8���;K{v1(J(���b��P�^���]�:��8�T��	��7�����|��誄o1Y������<}�A:���i�b�hU�,�Ś:'�vKȠNW���Ϻ��s8S2��o��@1F)�h*5� ��i6e^g�ɋIq�r��'���H[@_���c�6#]���@Y�T�J��e�#�	��&|�unS�#��;���Z�2_*$O2��%o�+�h��`~/4���&��N�H
�(�lYj���!H���aC����4�4��&R���7-6�]��Ƃ�e�v�9����-�)>|���m)�� ]�{�K��s����YN�4nH�Cm��$\�+>�0Z
Y���j#.���ke4�����$g����E��&��?5���׳I֡�G/c%?^���}�=��)
�߈��l}���lgL� ���`�	����PH"vKT�&��S��.��Ao�X���
��R9�s1MZEO5��Tw�!4Ց�ȗU�?#Q|m6}8V�r�[��r����Anq��MB�15SM�6]�/9th�V��+�v����՚᫭��q��F/�18�v� ������<��@�.�3�LLO�F쮊ss2<�sg�@�]�j���Q��Jp_�C�B�l��u/o�U]����1���L�)�����.q�y2C!�3�<K�F�)��-�)�����ݷ��K�~,��t��ì�H����A�$Z%��t�F���XԹ�t,v�G+������`�3����>��Y������%7���$�>���5�D9��q�ȯ�"���>�`�,�����HE�^autfj��x9e	�+B��ºb���!�w���뤥�"h�Fn�~y��A�>5�F��E���r��GaLmqSh�=C��P H�?�yɽ����q���wp,�S�b-d��@�Lٚ��E�\P3��L�-��"�����ǣx�����5`��O���lQ�W�X�� ��{��gC���.�0�W�@�]�q�F�)S���o�4\a�Y��� U	���
���'y�nF�v���Td������9zUsҡQ��E���<�q�*��Q�c�s�g�Ebc�,X���lS�OmT����/���;xO�bHN���8o�
� ��v����-
p�! kK+�s�;ԁ��A���ә'��]��{�3��o34-$u��f��k@��B">��2�uy��+Ҽ��hPHb������f�����3��в�5Ee���tm�������T��^�;1#f@^���3�� ��@8�\�^�w��!ʹ71�H0�c'~�4��ͼ���?ެHC7R��ډ���~"h;i>+X B�K�%hQb�ht�_�)��؃v��6|�i�V��{ԉa����aO4z���o��j�'S��5vA���)�)>��6p]����aZ
��y�6��J�V��c/����Kl��؈$X/24�H^с���72�FKk�*ĢrOw1n�ّ���R���Y�]�H%��%����e�)1g����a�VMH�NF��q�+7쌢�}�kT�cm|D¸Uk
+K;��au��Ķ�� ;�)��U�YO�	hw�,f/}��'��V�����O�o��Wu�%	�%&��%J{0wtXOO��H��i����ܘt��؆��9aW����*Ý�Y�4����=�<�����n MIǁ����:&��e�)�VS+���(
��T1�
c]�.W�s`�C�"��vY��h�m�5Y!�m�*a�,��r%�I<���TL����:ӯ��NN�zry�������*�{8���"��`�6@؎�J�n���aq��A����*8�rt�wbc�����:t�%tTp��8�M�k�#vC!�@Y�������x}�Gr��F���΄z��\����?I��I���+g�}��x���_͎d��F�b�󔣭��ϙ�����KG����a�L�Β�>0��J#���~f���-p�BH8��t��%8��K�� OQY���� <\���>!���^a�0w�(�����]�����v��\����o����RG��m��AUa�U�d��b����_� �SQG�\sB�	��؅K��PR�[2��3�R�w�H�X�`�h.	�o�h>�hkro��rg��\v��z��qd�����ܫ�h�bw&�Κq��L�o�|�֩�]O�v1��I��t�21`!���啬�g#�.�Tr�2��&����2Ӈ�S���2���s�4i1�W<�t)�b�hosjpJ�^�x��a\��?N~�9�;����%�wQ�&��1��9�2��Z���k�F�|B�v�ܪ�`��yd��tb�?�o �+&�#�?��j�-jcD׀,N��6�Թ���`L�0�F0��D��X��!n�c�I���]M���7�ؠA���k��T��}]�'3 ���B;Μ����!`|��<���[�õG>�}ʘ�uc��ݑ���j)�2��&X+�s��U�0�F�^lۖ����`;#�h�&%� ������`���,Qwm4x%a�L�qv� M�Vq`B�5�'�I�bg����ׯr�Z������A*'ֳ������˯9��������'ˏ{%��i���}��\zM�7-=ՌP����^��*����\���5�C}�Q-(�R@| v�ëN��6�&�.i{���=��@kgb.O�T���:�7��r�ݗ��Ջ�6M	\���Ch�A���P@���]^|�!���l��C�y�$��Yw�*�� K��p�G��O�&�[e��T��xpma��D�y�@��9��R8�Y��6�b{(�et�9��e�� ;9�j�dpUV�}�M8�����0����P|bv�U�k��B�>l$Sr�Wv}�s ���#Lvr䍊�&�j�h5霈֗����S�ԉ)�naU����['�O(Gv1YMnu9蛳F��x/㸌*��� �m�!���'-_��/�6їg����0TÜi��!�.c� �K�>�OP����,��0H�]��xuz}��\݇��`N۶�?R��z�[��P #�S˴��m�(��o���2�t�����'=U;] G1p@�����<Pb%?�c�;3���!̟��ϊU�9w����U�d|�_ټ[��Cb��2���?㰟B�V
8d����n���7ѡ�aO�-��b��8���MˠD�D�[x����_��<!���th�R���Գy�X�_U0.��,��e�������C��=������J�y�5Bk
�y��E���(�V6��?���|D��6=}�+�i�������=�SJ9��x�/�*Q����Jҝ��������c�6�@�פ	�YK�a6 �^�Qg#մ� 	�}�Ġ&�@t�شx�u.�L�Vl�V�����a �U⨹�G�:�e�ow��k9��� b4�z|�i='��E�(Yu��D셊ypK����*�:�!�]����v��n��+~IJ5�Q=�����;/��3�vM������+֘�j��ȳL�a�F��Ps.�Ÿ�duY.�X�QQq��B}(�H�.��<6*v��;����e���1�
k�|>{-��	{U��QBW��8�!lcd�5��Jh�a��c�;��D�"��d Ki��Ѷ�� �p]:-%O����V�$f������-3�8;��~J�n3Z��\�c5~pP�	�uR�����b��I�����a�А^���͏O��<y3c�v�H�Y�����d�+L;��dΝ�/�	V�[T�R|�B,��i���=�l>��"Z`[�HjV���W�>;a��>&���O�g�����$n��X�E��a�6:5DZ:kC7u�F��,��ٝ:i����t���
?���t�7T��4�BҥECf������.Y� G�5�����h�	�
7�H�
j&#Ov'{ �J�\?�b=�ڢQO�Rd�lЖ�J��y�v�ς�	G��0�nE���n���T�߫� ��5��o��ȞG�d�ɡ��������tw�}!��D���7Ń������Z���h��<���W�b��*��U&�ùb(����@��fA!�ކ�R,���j�	�nxѣ38K-F��o1���Ci�f�*rw�(y�/��q�t�����M`}�1ͩ%��pCИ����HM�ܻ��>���Hn��?���N�j�w�aDaiq�<�v�2����/���%,�y̙�[������CD|�rB|���6��u�&]�J��;r��
�r/#��2��g_��2 1���-oTѓ$*���b~����s��v�g�)�VB��PT����#�Ƴ7[?C��2	�Pڀ.u�u*�8�MC�v`��Ƿk��
�%�����z��#���#ŔĪ��)��I�F�h7d��z���!1�(�Y\��G�b֘&ؽ|��A�+�������aLSw��Qi��z�/����EU�$�u�g\��g�%����$�����(��k|�ѵ<�'����N�ћ�F�[�S�W��f-���N�g��h���X�ś�
5�/��;\>B�$ce�%��ef6�����\���K��|K�т�6�� ]٫�ִY�<�z �W��蓔�1�!��lf!y����?�9\rX��j�fQ,*6sM!�eV����9T��|��_�z僬s�<K��%�Vb�2���8�f���0 �ܝw���e� V�ڧ�^T�(�A�g$�f�f�/܂��qm�~�|u�b�ʀ8c����4��ߵvW�a�LQA���Q"��}Q'�K<�;�S$T�H�X�*�e(Gq���֌@O�u��o��#��
�b�W�+�,�dG�'�e��Q�sSwZ��u/��V1�����%�����Æ$y���*1��" �}7��ၞV���Dg߳��v:
�|�ב�f7�%�?�.�JUQ�YQ�0g(�r�M�b�P���Å��C�G?��#�vpz��:�V�����(t��������B�P�e�).��F6o��8� =�.N���ި��FI:2��[��c_TƦr
�=�|��;�/�r!`�i����*��©���x��<K�(m0+�Ǉ�s[Zm݋��#^�\VPp���A�.�DW�g�?a�+ ��{|��i��N�6fҩ���h{D��Y`1/湄�B�����z���4��e����6�#I�8qվP؃kp!4a*0����) ��L��*�����
Oݳ����� ݬoV�\���}BX���?Q#N�޼[�C{��s��N��a<tjJXR���a<Z�ډhD?�4���IG:d#=��L"�xT7xhb�1����zpU�yo�:�́��]�ƷPhO{ R��Ӿ�fڪ���,�Y�.KD���	��*Y�G��